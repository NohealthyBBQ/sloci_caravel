magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 302 316 336 394
rect 818 316 852 394
rect 1334 316 1368 394
rect 302 -500 336 -422
rect 818 -500 852 -422
rect 1334 -500 1368 -422
<< metal1 >>
rect 30 316 110 320
rect 30 264 44 316
rect 96 264 110 316
rect 30 260 110 264
rect 1050 316 1130 320
rect 1050 264 1064 316
rect 1116 264 1130 316
rect 1050 260 1130 264
rect 530 176 610 180
rect 530 124 544 176
rect 596 124 610 176
rect 530 120 610 124
rect 94 27 1318 73
rect 680 -133 740 27
rect 94 -180 1318 -133
rect 530 -224 610 -220
rect 530 -276 544 -224
rect 596 -276 610 -224
rect 530 -280 610 -276
rect 30 -364 110 -360
rect 30 -416 44 -364
rect 96 -416 110 -364
rect 30 -420 110 -416
rect 1050 -364 1130 -360
rect 1050 -416 1064 -364
rect 1116 -416 1130 -364
rect 1050 -420 1130 -416
<< via1 >>
rect 44 264 96 316
rect 1064 264 1116 316
rect 544 124 596 176
rect 544 -276 596 -224
rect 44 -416 96 -364
rect 1064 -416 1116 -364
<< metal2 >>
rect 40 320 100 330
rect 1060 320 1120 330
rect 40 316 1120 320
rect 40 264 44 316
rect 96 264 1064 316
rect 1116 264 1120 316
rect 40 260 1120 264
rect 40 250 100 260
rect 300 -220 360 260
rect 1060 250 1120 260
rect 540 180 600 190
rect 540 176 860 180
rect 540 124 544 176
rect 596 124 860 176
rect 540 120 860 124
rect 540 110 600 120
rect 540 -220 600 -210
rect 300 -224 600 -220
rect 300 -276 544 -224
rect 596 -276 600 -224
rect 300 -280 600 -276
rect 540 -290 600 -280
rect 40 -360 100 -350
rect 800 -360 860 120
rect 1060 -360 1120 -350
rect 40 -364 1120 -360
rect 40 -416 44 -364
rect 96 -416 1064 -364
rect 1116 -416 1120 -364
rect 40 -420 1120 -416
rect 40 -430 100 -420
rect 1060 -430 1120 -420
use sky130_fd_pr__pfet_01v8_lvt_MUVY4U  sky130_fd_pr__pfet_01v8_lvt_MUVY4U_0
timestamp 1663011646
transform 1 0 706 0 1 178
box -812 -284 812 284
use sky130_fd_pr__pfet_01v8_lvt_Q24T46  sky130_fd_pr__pfet_01v8_lvt_Q24T46_0
timestamp 1663011646
transform 1 0 706 0 1 -284
box -812 -284 812 284
<< end >>
