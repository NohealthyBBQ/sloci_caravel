magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal3 >>
rect -2150 3072 2149 3100
rect -2150 3008 2065 3072
rect 2129 3008 2149 3072
rect -2150 2992 2149 3008
rect -2150 2928 2065 2992
rect 2129 2928 2149 2992
rect -2150 2912 2149 2928
rect -2150 2848 2065 2912
rect 2129 2848 2149 2912
rect -2150 2832 2149 2848
rect -2150 2768 2065 2832
rect 2129 2768 2149 2832
rect -2150 2752 2149 2768
rect -2150 2688 2065 2752
rect 2129 2688 2149 2752
rect -2150 2672 2149 2688
rect -2150 2608 2065 2672
rect 2129 2608 2149 2672
rect -2150 2592 2149 2608
rect -2150 2528 2065 2592
rect 2129 2528 2149 2592
rect -2150 2512 2149 2528
rect -2150 2448 2065 2512
rect 2129 2448 2149 2512
rect -2150 2432 2149 2448
rect -2150 2368 2065 2432
rect 2129 2368 2149 2432
rect -2150 2352 2149 2368
rect -2150 2288 2065 2352
rect 2129 2288 2149 2352
rect -2150 2272 2149 2288
rect -2150 2208 2065 2272
rect 2129 2208 2149 2272
rect -2150 2192 2149 2208
rect -2150 2128 2065 2192
rect 2129 2128 2149 2192
rect -2150 2112 2149 2128
rect -2150 2048 2065 2112
rect 2129 2048 2149 2112
rect -2150 2032 2149 2048
rect -2150 1968 2065 2032
rect 2129 1968 2149 2032
rect -2150 1952 2149 1968
rect -2150 1888 2065 1952
rect 2129 1888 2149 1952
rect -2150 1872 2149 1888
rect -2150 1808 2065 1872
rect 2129 1808 2149 1872
rect -2150 1792 2149 1808
rect -2150 1728 2065 1792
rect 2129 1728 2149 1792
rect -2150 1712 2149 1728
rect -2150 1648 2065 1712
rect 2129 1648 2149 1712
rect -2150 1632 2149 1648
rect -2150 1568 2065 1632
rect 2129 1568 2149 1632
rect -2150 1552 2149 1568
rect -2150 1488 2065 1552
rect 2129 1488 2149 1552
rect -2150 1472 2149 1488
rect -2150 1408 2065 1472
rect 2129 1408 2149 1472
rect -2150 1392 2149 1408
rect -2150 1328 2065 1392
rect 2129 1328 2149 1392
rect -2150 1312 2149 1328
rect -2150 1248 2065 1312
rect 2129 1248 2149 1312
rect -2150 1232 2149 1248
rect -2150 1168 2065 1232
rect 2129 1168 2149 1232
rect -2150 1152 2149 1168
rect -2150 1088 2065 1152
rect 2129 1088 2149 1152
rect -2150 1072 2149 1088
rect -2150 1008 2065 1072
rect 2129 1008 2149 1072
rect -2150 992 2149 1008
rect -2150 928 2065 992
rect 2129 928 2149 992
rect -2150 912 2149 928
rect -2150 848 2065 912
rect 2129 848 2149 912
rect -2150 832 2149 848
rect -2150 768 2065 832
rect 2129 768 2149 832
rect -2150 752 2149 768
rect -2150 688 2065 752
rect 2129 688 2149 752
rect -2150 672 2149 688
rect -2150 608 2065 672
rect 2129 608 2149 672
rect -2150 592 2149 608
rect -2150 528 2065 592
rect 2129 528 2149 592
rect -2150 512 2149 528
rect -2150 448 2065 512
rect 2129 448 2149 512
rect -2150 432 2149 448
rect -2150 368 2065 432
rect 2129 368 2149 432
rect -2150 352 2149 368
rect -2150 288 2065 352
rect 2129 288 2149 352
rect -2150 272 2149 288
rect -2150 208 2065 272
rect 2129 208 2149 272
rect -2150 192 2149 208
rect -2150 128 2065 192
rect 2129 128 2149 192
rect -2150 112 2149 128
rect -2150 48 2065 112
rect 2129 48 2149 112
rect -2150 32 2149 48
rect -2150 -32 2065 32
rect 2129 -32 2149 32
rect -2150 -48 2149 -32
rect -2150 -112 2065 -48
rect 2129 -112 2149 -48
rect -2150 -128 2149 -112
rect -2150 -192 2065 -128
rect 2129 -192 2149 -128
rect -2150 -208 2149 -192
rect -2150 -272 2065 -208
rect 2129 -272 2149 -208
rect -2150 -288 2149 -272
rect -2150 -352 2065 -288
rect 2129 -352 2149 -288
rect -2150 -368 2149 -352
rect -2150 -432 2065 -368
rect 2129 -432 2149 -368
rect -2150 -448 2149 -432
rect -2150 -512 2065 -448
rect 2129 -512 2149 -448
rect -2150 -528 2149 -512
rect -2150 -592 2065 -528
rect 2129 -592 2149 -528
rect -2150 -608 2149 -592
rect -2150 -672 2065 -608
rect 2129 -672 2149 -608
rect -2150 -688 2149 -672
rect -2150 -752 2065 -688
rect 2129 -752 2149 -688
rect -2150 -768 2149 -752
rect -2150 -832 2065 -768
rect 2129 -832 2149 -768
rect -2150 -848 2149 -832
rect -2150 -912 2065 -848
rect 2129 -912 2149 -848
rect -2150 -928 2149 -912
rect -2150 -992 2065 -928
rect 2129 -992 2149 -928
rect -2150 -1008 2149 -992
rect -2150 -1072 2065 -1008
rect 2129 -1072 2149 -1008
rect -2150 -1088 2149 -1072
rect -2150 -1152 2065 -1088
rect 2129 -1152 2149 -1088
rect -2150 -1168 2149 -1152
rect -2150 -1232 2065 -1168
rect 2129 -1232 2149 -1168
rect -2150 -1248 2149 -1232
rect -2150 -1312 2065 -1248
rect 2129 -1312 2149 -1248
rect -2150 -1328 2149 -1312
rect -2150 -1392 2065 -1328
rect 2129 -1392 2149 -1328
rect -2150 -1408 2149 -1392
rect -2150 -1472 2065 -1408
rect 2129 -1472 2149 -1408
rect -2150 -1488 2149 -1472
rect -2150 -1552 2065 -1488
rect 2129 -1552 2149 -1488
rect -2150 -1568 2149 -1552
rect -2150 -1632 2065 -1568
rect 2129 -1632 2149 -1568
rect -2150 -1648 2149 -1632
rect -2150 -1712 2065 -1648
rect 2129 -1712 2149 -1648
rect -2150 -1728 2149 -1712
rect -2150 -1792 2065 -1728
rect 2129 -1792 2149 -1728
rect -2150 -1808 2149 -1792
rect -2150 -1872 2065 -1808
rect 2129 -1872 2149 -1808
rect -2150 -1888 2149 -1872
rect -2150 -1952 2065 -1888
rect 2129 -1952 2149 -1888
rect -2150 -1968 2149 -1952
rect -2150 -2032 2065 -1968
rect 2129 -2032 2149 -1968
rect -2150 -2048 2149 -2032
rect -2150 -2112 2065 -2048
rect 2129 -2112 2149 -2048
rect -2150 -2128 2149 -2112
rect -2150 -2192 2065 -2128
rect 2129 -2192 2149 -2128
rect -2150 -2208 2149 -2192
rect -2150 -2272 2065 -2208
rect 2129 -2272 2149 -2208
rect -2150 -2288 2149 -2272
rect -2150 -2352 2065 -2288
rect 2129 -2352 2149 -2288
rect -2150 -2368 2149 -2352
rect -2150 -2432 2065 -2368
rect 2129 -2432 2149 -2368
rect -2150 -2448 2149 -2432
rect -2150 -2512 2065 -2448
rect 2129 -2512 2149 -2448
rect -2150 -2528 2149 -2512
rect -2150 -2592 2065 -2528
rect 2129 -2592 2149 -2528
rect -2150 -2608 2149 -2592
rect -2150 -2672 2065 -2608
rect 2129 -2672 2149 -2608
rect -2150 -2688 2149 -2672
rect -2150 -2752 2065 -2688
rect 2129 -2752 2149 -2688
rect -2150 -2768 2149 -2752
rect -2150 -2832 2065 -2768
rect 2129 -2832 2149 -2768
rect -2150 -2848 2149 -2832
rect -2150 -2912 2065 -2848
rect 2129 -2912 2149 -2848
rect -2150 -2928 2149 -2912
rect -2150 -2992 2065 -2928
rect 2129 -2992 2149 -2928
rect -2150 -3008 2149 -2992
rect -2150 -3072 2065 -3008
rect 2129 -3072 2149 -3008
rect -2150 -3100 2149 -3072
<< via3 >>
rect 2065 3008 2129 3072
rect 2065 2928 2129 2992
rect 2065 2848 2129 2912
rect 2065 2768 2129 2832
rect 2065 2688 2129 2752
rect 2065 2608 2129 2672
rect 2065 2528 2129 2592
rect 2065 2448 2129 2512
rect 2065 2368 2129 2432
rect 2065 2288 2129 2352
rect 2065 2208 2129 2272
rect 2065 2128 2129 2192
rect 2065 2048 2129 2112
rect 2065 1968 2129 2032
rect 2065 1888 2129 1952
rect 2065 1808 2129 1872
rect 2065 1728 2129 1792
rect 2065 1648 2129 1712
rect 2065 1568 2129 1632
rect 2065 1488 2129 1552
rect 2065 1408 2129 1472
rect 2065 1328 2129 1392
rect 2065 1248 2129 1312
rect 2065 1168 2129 1232
rect 2065 1088 2129 1152
rect 2065 1008 2129 1072
rect 2065 928 2129 992
rect 2065 848 2129 912
rect 2065 768 2129 832
rect 2065 688 2129 752
rect 2065 608 2129 672
rect 2065 528 2129 592
rect 2065 448 2129 512
rect 2065 368 2129 432
rect 2065 288 2129 352
rect 2065 208 2129 272
rect 2065 128 2129 192
rect 2065 48 2129 112
rect 2065 -32 2129 32
rect 2065 -112 2129 -48
rect 2065 -192 2129 -128
rect 2065 -272 2129 -208
rect 2065 -352 2129 -288
rect 2065 -432 2129 -368
rect 2065 -512 2129 -448
rect 2065 -592 2129 -528
rect 2065 -672 2129 -608
rect 2065 -752 2129 -688
rect 2065 -832 2129 -768
rect 2065 -912 2129 -848
rect 2065 -992 2129 -928
rect 2065 -1072 2129 -1008
rect 2065 -1152 2129 -1088
rect 2065 -1232 2129 -1168
rect 2065 -1312 2129 -1248
rect 2065 -1392 2129 -1328
rect 2065 -1472 2129 -1408
rect 2065 -1552 2129 -1488
rect 2065 -1632 2129 -1568
rect 2065 -1712 2129 -1648
rect 2065 -1792 2129 -1728
rect 2065 -1872 2129 -1808
rect 2065 -1952 2129 -1888
rect 2065 -2032 2129 -1968
rect 2065 -2112 2129 -2048
rect 2065 -2192 2129 -2128
rect 2065 -2272 2129 -2208
rect 2065 -2352 2129 -2288
rect 2065 -2432 2129 -2368
rect 2065 -2512 2129 -2448
rect 2065 -2592 2129 -2528
rect 2065 -2672 2129 -2608
rect 2065 -2752 2129 -2688
rect 2065 -2832 2129 -2768
rect 2065 -2912 2129 -2848
rect 2065 -2992 2129 -2928
rect 2065 -3072 2129 -3008
<< mimcap >>
rect -2050 2952 1950 3000
rect -2050 -2952 -2002 2952
rect 1902 -2952 1950 2952
rect -2050 -3000 1950 -2952
<< mimcapcontact >>
rect -2002 -2952 1902 2952
<< metal4 >>
rect 2049 3072 2145 3088
rect 2049 3008 2065 3072
rect 2129 3008 2145 3072
rect 2049 2992 2145 3008
rect -2011 2952 1911 2961
rect -2011 -2952 -2002 2952
rect 1902 -2952 1911 2952
rect -2011 -2961 1911 -2952
rect 2049 2928 2065 2992
rect 2129 2928 2145 2992
rect 2049 2912 2145 2928
rect 2049 2848 2065 2912
rect 2129 2848 2145 2912
rect 2049 2832 2145 2848
rect 2049 2768 2065 2832
rect 2129 2768 2145 2832
rect 2049 2752 2145 2768
rect 2049 2688 2065 2752
rect 2129 2688 2145 2752
rect 2049 2672 2145 2688
rect 2049 2608 2065 2672
rect 2129 2608 2145 2672
rect 2049 2592 2145 2608
rect 2049 2528 2065 2592
rect 2129 2528 2145 2592
rect 2049 2512 2145 2528
rect 2049 2448 2065 2512
rect 2129 2448 2145 2512
rect 2049 2432 2145 2448
rect 2049 2368 2065 2432
rect 2129 2368 2145 2432
rect 2049 2352 2145 2368
rect 2049 2288 2065 2352
rect 2129 2288 2145 2352
rect 2049 2272 2145 2288
rect 2049 2208 2065 2272
rect 2129 2208 2145 2272
rect 2049 2192 2145 2208
rect 2049 2128 2065 2192
rect 2129 2128 2145 2192
rect 2049 2112 2145 2128
rect 2049 2048 2065 2112
rect 2129 2048 2145 2112
rect 2049 2032 2145 2048
rect 2049 1968 2065 2032
rect 2129 1968 2145 2032
rect 2049 1952 2145 1968
rect 2049 1888 2065 1952
rect 2129 1888 2145 1952
rect 2049 1872 2145 1888
rect 2049 1808 2065 1872
rect 2129 1808 2145 1872
rect 2049 1792 2145 1808
rect 2049 1728 2065 1792
rect 2129 1728 2145 1792
rect 2049 1712 2145 1728
rect 2049 1648 2065 1712
rect 2129 1648 2145 1712
rect 2049 1632 2145 1648
rect 2049 1568 2065 1632
rect 2129 1568 2145 1632
rect 2049 1552 2145 1568
rect 2049 1488 2065 1552
rect 2129 1488 2145 1552
rect 2049 1472 2145 1488
rect 2049 1408 2065 1472
rect 2129 1408 2145 1472
rect 2049 1392 2145 1408
rect 2049 1328 2065 1392
rect 2129 1328 2145 1392
rect 2049 1312 2145 1328
rect 2049 1248 2065 1312
rect 2129 1248 2145 1312
rect 2049 1232 2145 1248
rect 2049 1168 2065 1232
rect 2129 1168 2145 1232
rect 2049 1152 2145 1168
rect 2049 1088 2065 1152
rect 2129 1088 2145 1152
rect 2049 1072 2145 1088
rect 2049 1008 2065 1072
rect 2129 1008 2145 1072
rect 2049 992 2145 1008
rect 2049 928 2065 992
rect 2129 928 2145 992
rect 2049 912 2145 928
rect 2049 848 2065 912
rect 2129 848 2145 912
rect 2049 832 2145 848
rect 2049 768 2065 832
rect 2129 768 2145 832
rect 2049 752 2145 768
rect 2049 688 2065 752
rect 2129 688 2145 752
rect 2049 672 2145 688
rect 2049 608 2065 672
rect 2129 608 2145 672
rect 2049 592 2145 608
rect 2049 528 2065 592
rect 2129 528 2145 592
rect 2049 512 2145 528
rect 2049 448 2065 512
rect 2129 448 2145 512
rect 2049 432 2145 448
rect 2049 368 2065 432
rect 2129 368 2145 432
rect 2049 352 2145 368
rect 2049 288 2065 352
rect 2129 288 2145 352
rect 2049 272 2145 288
rect 2049 208 2065 272
rect 2129 208 2145 272
rect 2049 192 2145 208
rect 2049 128 2065 192
rect 2129 128 2145 192
rect 2049 112 2145 128
rect 2049 48 2065 112
rect 2129 48 2145 112
rect 2049 32 2145 48
rect 2049 -32 2065 32
rect 2129 -32 2145 32
rect 2049 -48 2145 -32
rect 2049 -112 2065 -48
rect 2129 -112 2145 -48
rect 2049 -128 2145 -112
rect 2049 -192 2065 -128
rect 2129 -192 2145 -128
rect 2049 -208 2145 -192
rect 2049 -272 2065 -208
rect 2129 -272 2145 -208
rect 2049 -288 2145 -272
rect 2049 -352 2065 -288
rect 2129 -352 2145 -288
rect 2049 -368 2145 -352
rect 2049 -432 2065 -368
rect 2129 -432 2145 -368
rect 2049 -448 2145 -432
rect 2049 -512 2065 -448
rect 2129 -512 2145 -448
rect 2049 -528 2145 -512
rect 2049 -592 2065 -528
rect 2129 -592 2145 -528
rect 2049 -608 2145 -592
rect 2049 -672 2065 -608
rect 2129 -672 2145 -608
rect 2049 -688 2145 -672
rect 2049 -752 2065 -688
rect 2129 -752 2145 -688
rect 2049 -768 2145 -752
rect 2049 -832 2065 -768
rect 2129 -832 2145 -768
rect 2049 -848 2145 -832
rect 2049 -912 2065 -848
rect 2129 -912 2145 -848
rect 2049 -928 2145 -912
rect 2049 -992 2065 -928
rect 2129 -992 2145 -928
rect 2049 -1008 2145 -992
rect 2049 -1072 2065 -1008
rect 2129 -1072 2145 -1008
rect 2049 -1088 2145 -1072
rect 2049 -1152 2065 -1088
rect 2129 -1152 2145 -1088
rect 2049 -1168 2145 -1152
rect 2049 -1232 2065 -1168
rect 2129 -1232 2145 -1168
rect 2049 -1248 2145 -1232
rect 2049 -1312 2065 -1248
rect 2129 -1312 2145 -1248
rect 2049 -1328 2145 -1312
rect 2049 -1392 2065 -1328
rect 2129 -1392 2145 -1328
rect 2049 -1408 2145 -1392
rect 2049 -1472 2065 -1408
rect 2129 -1472 2145 -1408
rect 2049 -1488 2145 -1472
rect 2049 -1552 2065 -1488
rect 2129 -1552 2145 -1488
rect 2049 -1568 2145 -1552
rect 2049 -1632 2065 -1568
rect 2129 -1632 2145 -1568
rect 2049 -1648 2145 -1632
rect 2049 -1712 2065 -1648
rect 2129 -1712 2145 -1648
rect 2049 -1728 2145 -1712
rect 2049 -1792 2065 -1728
rect 2129 -1792 2145 -1728
rect 2049 -1808 2145 -1792
rect 2049 -1872 2065 -1808
rect 2129 -1872 2145 -1808
rect 2049 -1888 2145 -1872
rect 2049 -1952 2065 -1888
rect 2129 -1952 2145 -1888
rect 2049 -1968 2145 -1952
rect 2049 -2032 2065 -1968
rect 2129 -2032 2145 -1968
rect 2049 -2048 2145 -2032
rect 2049 -2112 2065 -2048
rect 2129 -2112 2145 -2048
rect 2049 -2128 2145 -2112
rect 2049 -2192 2065 -2128
rect 2129 -2192 2145 -2128
rect 2049 -2208 2145 -2192
rect 2049 -2272 2065 -2208
rect 2129 -2272 2145 -2208
rect 2049 -2288 2145 -2272
rect 2049 -2352 2065 -2288
rect 2129 -2352 2145 -2288
rect 2049 -2368 2145 -2352
rect 2049 -2432 2065 -2368
rect 2129 -2432 2145 -2368
rect 2049 -2448 2145 -2432
rect 2049 -2512 2065 -2448
rect 2129 -2512 2145 -2448
rect 2049 -2528 2145 -2512
rect 2049 -2592 2065 -2528
rect 2129 -2592 2145 -2528
rect 2049 -2608 2145 -2592
rect 2049 -2672 2065 -2608
rect 2129 -2672 2145 -2608
rect 2049 -2688 2145 -2672
rect 2049 -2752 2065 -2688
rect 2129 -2752 2145 -2688
rect 2049 -2768 2145 -2752
rect 2049 -2832 2065 -2768
rect 2129 -2832 2145 -2768
rect 2049 -2848 2145 -2832
rect 2049 -2912 2065 -2848
rect 2129 -2912 2145 -2848
rect 2049 -2928 2145 -2912
rect 2049 -2992 2065 -2928
rect 2129 -2992 2145 -2928
rect 2049 -3008 2145 -2992
rect 2049 -3072 2065 -3008
rect 2129 -3072 2145 -3008
rect 2049 -3088 2145 -3072
<< properties >>
string FIXED_BBOX -2150 -3100 2050 3100
<< end >>
