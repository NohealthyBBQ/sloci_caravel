magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect 17100 7240 19040 7245
rect 17710 5070 19040 7240
rect 17710 4990 17780 5070
rect 18360 4990 18420 5070
rect 18620 5020 19040 5070
rect 19035 4990 19040 5020
rect 18180 4384 18600 4390
rect 17930 210 18350 4384
rect 20550 2400 20750 5650
<< locali >>
rect 17670 7175 17825 7215
rect 18315 7170 18470 7210
rect 18970 6975 20025 7020
rect 19990 6180 20025 6975
rect 20520 5545 20775 5580
rect 17535 4310 17570 5060
rect 17670 5030 17825 5070
rect 18070 4350 18105 5060
rect 18185 4350 18220 5060
rect 18320 5030 18475 5070
rect 18070 4315 18220 4350
rect 18715 4315 18750 5065
rect 18185 4310 18220 4315
rect 19075 4105 19110 4270
rect 19870 4105 19905 4270
rect 20735 4070 20770 4075
rect 19985 3930 20020 4070
rect 20515 4035 20775 4070
rect 20520 3980 20555 4035
rect 20735 3980 20770 4035
rect 20510 3935 20770 3980
rect 21265 3940 21300 4080
rect 20515 2435 20770 2470
rect 18070 245 18220 280
rect 18070 -100 18220 -65
rect 19070 -100 19115 790
rect 19370 -95 19410 780
rect 18070 -615 18220 -580
<< metal1 >>
rect 17220 7150 20470 7220
rect 17220 5180 17280 7150
rect 17310 7106 17400 7120
rect 17310 7054 17329 7106
rect 17381 7100 17400 7106
rect 17381 7054 17530 7100
rect 17310 7050 17530 7054
rect 17310 7040 17400 7050
rect 17440 6976 17530 6990
rect 17440 6970 17459 6976
rect 17310 6924 17459 6970
rect 17511 6924 17530 6976
rect 17310 6920 17530 6924
rect 17440 6910 17530 6920
rect 17310 6846 17400 6860
rect 17310 6794 17329 6846
rect 17381 6840 17400 6846
rect 17381 6794 17530 6840
rect 17310 6790 17530 6794
rect 17310 6780 17400 6790
rect 17440 6720 17530 6730
rect 17310 6716 17530 6720
rect 17310 6670 17459 6716
rect 17440 6664 17459 6670
rect 17511 6664 17530 6716
rect 17440 6650 17530 6664
rect 17310 6590 17400 6600
rect 17310 6586 17530 6590
rect 17310 6534 17329 6586
rect 17381 6540 17530 6586
rect 17381 6534 17400 6540
rect 17310 6520 17400 6534
rect 17440 6460 17530 6470
rect 17310 6456 17530 6460
rect 17310 6410 17459 6456
rect 17440 6404 17459 6410
rect 17511 6404 17530 6456
rect 17440 6390 17530 6404
rect 17310 6330 17400 6340
rect 17310 6326 17530 6330
rect 17310 6274 17329 6326
rect 17381 6280 17530 6326
rect 17381 6274 17400 6280
rect 17310 6260 17400 6274
rect 17440 6206 17530 6220
rect 17440 6200 17459 6206
rect 17310 6160 17459 6200
rect 17440 6154 17459 6160
rect 17511 6154 17530 6206
rect 17440 6140 17530 6154
rect 17310 6080 17400 6090
rect 17310 6076 17530 6080
rect 17310 6024 17329 6076
rect 17381 6030 17530 6076
rect 17381 6024 17400 6030
rect 17310 6010 17400 6024
rect 17440 5956 17530 5970
rect 17440 5950 17459 5956
rect 17310 5904 17459 5950
rect 17511 5904 17530 5956
rect 17310 5900 17530 5904
rect 17440 5890 17530 5900
rect 17310 5826 17400 5840
rect 17310 5774 17329 5826
rect 17381 5820 17400 5826
rect 17381 5774 17530 5820
rect 17310 5770 17530 5774
rect 17310 5760 17400 5770
rect 17440 5696 17530 5710
rect 17440 5690 17459 5696
rect 17310 5644 17459 5690
rect 17511 5644 17530 5696
rect 17310 5640 17530 5644
rect 17440 5630 17530 5640
rect 17310 5566 17400 5580
rect 17310 5514 17329 5566
rect 17381 5560 17400 5566
rect 17381 5520 17530 5560
rect 17381 5514 17400 5520
rect 17310 5500 17400 5514
rect 17440 5440 17530 5450
rect 17310 5436 17530 5440
rect 17310 5390 17459 5436
rect 17440 5384 17459 5390
rect 17511 5384 17530 5436
rect 17440 5370 17530 5384
rect 17310 5310 17400 5320
rect 17310 5306 17530 5310
rect 17310 5254 17329 5306
rect 17381 5260 17530 5306
rect 17381 5254 17400 5260
rect 17310 5240 17400 5254
rect 17440 5180 17530 5190
rect 17560 5180 17620 7150
rect 17870 5180 17930 7150
rect 17960 7106 18050 7120
rect 17960 7054 17979 7106
rect 18031 7100 18050 7106
rect 18031 7054 18180 7100
rect 17960 7050 18180 7054
rect 17960 7040 18050 7050
rect 18090 6976 18180 6990
rect 18090 6972 18109 6976
rect 17969 6970 18109 6972
rect 17960 6924 18109 6970
rect 18161 6924 18180 6976
rect 17960 6920 18180 6924
rect 18090 6910 18180 6920
rect 17960 6846 18050 6860
rect 17960 6794 17979 6846
rect 18031 6844 18050 6846
rect 18031 6840 18169 6844
rect 18031 6794 18180 6840
rect 17960 6790 18180 6794
rect 17960 6780 18050 6790
rect 18090 6720 18180 6730
rect 17960 6716 18180 6720
rect 17960 6670 18109 6716
rect 18090 6664 18109 6670
rect 18161 6664 18180 6716
rect 18090 6650 18180 6664
rect 17960 6590 18050 6600
rect 17960 6586 18180 6590
rect 17960 6534 17979 6586
rect 18031 6540 18180 6586
rect 18031 6534 18050 6540
rect 17960 6520 18050 6534
rect 18090 6460 18180 6470
rect 17960 6456 18180 6460
rect 17960 6410 18109 6456
rect 18090 6404 18109 6410
rect 18161 6404 18180 6456
rect 18090 6390 18180 6404
rect 17960 6332 18050 6340
rect 17960 6330 18169 6332
rect 17960 6326 18180 6330
rect 17960 6274 17979 6326
rect 18031 6280 18180 6326
rect 18031 6274 18050 6280
rect 17960 6260 18050 6274
rect 18090 6206 18180 6220
rect 18090 6204 18109 6206
rect 17969 6200 18109 6204
rect 17960 6160 18109 6200
rect 17969 6158 18109 6160
rect 18090 6154 18109 6158
rect 18161 6154 18180 6206
rect 18090 6140 18180 6154
rect 17960 6080 18050 6090
rect 17960 6076 18180 6080
rect 17960 6024 17979 6076
rect 18031 6030 18180 6076
rect 18031 6024 18050 6030
rect 17960 6010 18050 6024
rect 18090 5956 18180 5970
rect 18090 5950 18109 5956
rect 17960 5904 18109 5950
rect 18161 5904 18180 5956
rect 17960 5900 18180 5904
rect 18090 5890 18180 5900
rect 17960 5826 18050 5840
rect 17960 5774 17979 5826
rect 18031 5820 18050 5826
rect 18031 5774 18180 5820
rect 17960 5770 18180 5774
rect 17960 5760 18050 5770
rect 18090 5696 18180 5710
rect 18090 5692 18109 5696
rect 17969 5690 18109 5692
rect 17960 5644 18109 5690
rect 18161 5644 18180 5696
rect 17960 5640 18180 5644
rect 18090 5630 18180 5640
rect 17960 5566 18050 5580
rect 17960 5514 17979 5566
rect 18031 5564 18050 5566
rect 18031 5560 18169 5564
rect 18031 5520 18180 5560
rect 18031 5518 18169 5520
rect 18031 5514 18050 5518
rect 17960 5500 18050 5514
rect 18090 5440 18180 5450
rect 17960 5436 18180 5440
rect 17960 5390 18109 5436
rect 18090 5384 18109 5390
rect 18161 5384 18180 5436
rect 18090 5370 18180 5384
rect 17960 5310 18050 5320
rect 17960 5306 18180 5310
rect 17960 5254 17979 5306
rect 18031 5260 18180 5306
rect 18031 5254 18050 5260
rect 17960 5240 18050 5254
rect 18090 5180 18180 5190
rect 18210 5180 18270 7150
rect 18520 5180 18580 7150
rect 18610 7106 18700 7120
rect 18610 7054 18629 7106
rect 18681 7100 18700 7106
rect 18681 7054 18830 7100
rect 18610 7050 18830 7054
rect 18610 7040 18700 7050
rect 18740 6976 18830 6990
rect 18740 6972 18759 6976
rect 18619 6970 18759 6972
rect 18610 6924 18759 6970
rect 18811 6924 18830 6976
rect 18610 6920 18830 6924
rect 18740 6910 18830 6920
rect 18610 6846 18700 6860
rect 18610 6794 18629 6846
rect 18681 6844 18700 6846
rect 18681 6840 18819 6844
rect 18681 6794 18830 6840
rect 18610 6790 18830 6794
rect 18610 6780 18700 6790
rect 18740 6720 18830 6730
rect 18610 6716 18830 6720
rect 18610 6670 18759 6716
rect 18740 6664 18759 6670
rect 18811 6664 18830 6716
rect 18740 6650 18830 6664
rect 18610 6590 18700 6600
rect 18610 6586 18830 6590
rect 18610 6534 18629 6586
rect 18681 6540 18830 6586
rect 18681 6534 18700 6540
rect 18610 6520 18700 6534
rect 18740 6460 18830 6470
rect 18610 6456 18830 6460
rect 18610 6410 18759 6456
rect 18740 6404 18759 6410
rect 18811 6404 18830 6456
rect 18740 6390 18830 6404
rect 18610 6332 18700 6340
rect 18610 6330 18819 6332
rect 18610 6326 18830 6330
rect 18610 6274 18629 6326
rect 18681 6280 18830 6326
rect 18681 6274 18700 6280
rect 18610 6260 18700 6274
rect 18740 6206 18830 6220
rect 18740 6204 18759 6206
rect 18619 6200 18759 6204
rect 18610 6160 18759 6200
rect 18619 6158 18759 6160
rect 18740 6154 18759 6158
rect 18811 6154 18830 6206
rect 18740 6140 18830 6154
rect 18610 6080 18700 6090
rect 18610 6076 18830 6080
rect 18610 6024 18629 6076
rect 18681 6030 18830 6076
rect 18681 6024 18700 6030
rect 18610 6010 18700 6024
rect 18740 5956 18830 5970
rect 18740 5950 18759 5956
rect 18610 5904 18759 5950
rect 18811 5904 18830 5956
rect 18610 5900 18830 5904
rect 18740 5890 18830 5900
rect 18610 5826 18700 5840
rect 18610 5774 18629 5826
rect 18681 5820 18700 5826
rect 18681 5774 18830 5820
rect 18610 5770 18830 5774
rect 18610 5760 18700 5770
rect 18740 5696 18830 5710
rect 18740 5692 18759 5696
rect 18619 5690 18759 5692
rect 18610 5644 18759 5690
rect 18811 5644 18830 5696
rect 18610 5640 18830 5644
rect 18740 5630 18830 5640
rect 18610 5566 18700 5580
rect 18610 5514 18629 5566
rect 18681 5564 18700 5566
rect 18681 5560 18819 5564
rect 18681 5520 18830 5560
rect 18681 5518 18819 5520
rect 18681 5514 18700 5518
rect 18610 5500 18700 5514
rect 18740 5440 18830 5450
rect 18610 5436 18830 5440
rect 18610 5390 18759 5436
rect 18740 5384 18759 5390
rect 18811 5384 18830 5436
rect 18740 5370 18830 5384
rect 18610 5310 18700 5320
rect 18610 5306 18830 5310
rect 18610 5254 18629 5306
rect 18681 5260 18830 5306
rect 18681 5254 18700 5260
rect 18610 5240 18700 5254
rect 18740 5180 18830 5190
rect 18860 5180 18920 7150
rect 19235 6703 19740 6710
rect 19235 6331 19237 6703
rect 19737 6331 19740 6703
rect 19235 6325 19740 6331
rect 20410 6220 20470 7150
rect 20070 6160 20470 6220
rect 17310 5176 17530 5180
rect 17310 5130 17459 5176
rect 17440 5124 17459 5130
rect 17511 5124 17530 5176
rect 17960 5176 18180 5180
rect 17960 5130 18109 5176
rect 17440 5110 17530 5124
rect 18090 5124 18109 5130
rect 18161 5124 18180 5176
rect 18610 5176 18830 5180
rect 18610 5130 18759 5176
rect 18090 5110 18180 5124
rect 18740 5124 18759 5130
rect 18811 5124 18830 5176
rect 18740 5110 18830 5124
rect 17100 4310 18020 4370
rect 17620 400 17680 4310
rect 17710 4241 17790 4260
rect 17710 4189 17724 4241
rect 17776 4189 17790 4241
rect 17860 4190 17930 4240
rect 17710 4170 17790 4189
rect 17850 4111 17930 4130
rect 17850 4110 17864 4111
rect 17710 4060 17864 4110
rect 17850 4059 17864 4060
rect 17916 4059 17930 4111
rect 17850 4040 17930 4059
rect 17710 3990 17790 4000
rect 17710 3981 17930 3990
rect 17710 3929 17724 3981
rect 17776 3940 17930 3981
rect 17776 3929 17790 3940
rect 17710 3910 17790 3929
rect 17850 3861 17930 3880
rect 17850 3860 17864 3861
rect 17710 3810 17864 3860
rect 17850 3809 17864 3810
rect 17916 3809 17930 3861
rect 17850 3790 17930 3809
rect 17710 3731 17790 3750
rect 17710 3679 17724 3731
rect 17776 3730 17790 3731
rect 17776 3680 17930 3730
rect 17776 3679 17790 3680
rect 17710 3660 17790 3679
rect 17850 3601 17930 3620
rect 17850 3600 17864 3601
rect 17710 3550 17864 3600
rect 17850 3549 17864 3550
rect 17916 3549 17930 3601
rect 17850 3530 17930 3549
rect 17710 3471 17790 3490
rect 17710 3419 17724 3471
rect 17776 3470 17790 3471
rect 17776 3420 17930 3470
rect 17776 3419 17790 3420
rect 17710 3400 17790 3419
rect 17850 3351 17930 3370
rect 17850 3350 17864 3351
rect 17710 3300 17864 3350
rect 17850 3299 17864 3300
rect 17916 3299 17930 3351
rect 17850 3280 17930 3299
rect 17710 3221 17790 3240
rect 17710 3169 17724 3221
rect 17776 3220 17790 3221
rect 17776 3170 17930 3220
rect 17776 3169 17790 3170
rect 17710 3150 17790 3169
rect 17850 3091 17930 3110
rect 17850 3090 17864 3091
rect 17710 3040 17864 3090
rect 17850 3039 17864 3040
rect 17916 3039 17930 3091
rect 17850 3020 17930 3039
rect 17710 2961 17790 2980
rect 17710 2909 17724 2961
rect 17776 2960 17790 2961
rect 17776 2910 17930 2960
rect 17776 2909 17790 2910
rect 17710 2890 17790 2909
rect 17850 2831 17930 2850
rect 17850 2830 17864 2831
rect 17710 2780 17864 2830
rect 17850 2779 17864 2780
rect 17916 2779 17930 2831
rect 17850 2760 17930 2779
rect 17710 2711 17790 2730
rect 17710 2659 17724 2711
rect 17776 2710 17790 2711
rect 17776 2659 17930 2710
rect 17710 2650 17930 2659
rect 17710 2640 17790 2650
rect 17850 2581 17930 2600
rect 17850 2580 17864 2581
rect 17710 2530 17864 2580
rect 17850 2529 17864 2530
rect 17916 2529 17930 2581
rect 17850 2510 17930 2529
rect 17710 2451 17790 2470
rect 17710 2399 17724 2451
rect 17776 2450 17790 2451
rect 17776 2400 17930 2450
rect 17776 2399 17790 2400
rect 17710 2380 17790 2399
rect 17850 2321 17930 2340
rect 17850 2320 17864 2321
rect 17710 2270 17864 2320
rect 17850 2269 17864 2270
rect 17916 2269 17930 2321
rect 17850 2250 17930 2269
rect 17710 2200 17790 2210
rect 17710 2191 17930 2200
rect 17710 2139 17724 2191
rect 17776 2140 17930 2191
rect 17776 2139 17790 2140
rect 17710 2120 17790 2139
rect 17850 2071 17930 2090
rect 17850 2070 17864 2071
rect 17710 2019 17864 2070
rect 17916 2019 17930 2071
rect 17710 2010 17930 2019
rect 17850 2000 17930 2010
rect 17710 1941 17790 1960
rect 17710 1889 17724 1941
rect 17776 1940 17790 1941
rect 17776 1890 17930 1940
rect 17776 1889 17790 1890
rect 17710 1870 17790 1889
rect 17850 1811 17930 1830
rect 17850 1810 17864 1811
rect 17710 1760 17864 1810
rect 17850 1759 17864 1760
rect 17916 1759 17930 1811
rect 17850 1740 17930 1759
rect 17710 1681 17790 1700
rect 17710 1629 17724 1681
rect 17776 1680 17790 1681
rect 17776 1630 17930 1680
rect 17776 1629 17790 1630
rect 17710 1610 17790 1629
rect 17850 1551 17930 1570
rect 17850 1550 17864 1551
rect 17710 1510 17864 1550
rect 17850 1499 17864 1510
rect 17916 1499 17930 1551
rect 17850 1480 17930 1499
rect 17710 1430 17790 1440
rect 17710 1421 17930 1430
rect 17710 1369 17724 1421
rect 17776 1380 17930 1421
rect 17776 1369 17790 1380
rect 17710 1350 17790 1369
rect 17850 1301 17930 1320
rect 17850 1300 17864 1301
rect 17710 1250 17864 1300
rect 17850 1249 17864 1250
rect 17916 1249 17930 1301
rect 17850 1230 17930 1249
rect 17710 1171 17790 1190
rect 17710 1119 17724 1171
rect 17776 1170 17790 1171
rect 17776 1120 17930 1170
rect 17776 1119 17790 1120
rect 17710 1100 17790 1119
rect 17850 1041 17930 1060
rect 17850 1040 17864 1041
rect 17710 990 17864 1040
rect 17850 989 17864 990
rect 17916 989 17930 1041
rect 17850 970 17930 989
rect 17710 911 17790 930
rect 17710 859 17724 911
rect 17776 910 17790 911
rect 17776 860 17930 910
rect 17776 859 17790 860
rect 17710 840 17790 859
rect 17850 791 17930 810
rect 17850 790 17864 791
rect 17710 739 17864 790
rect 17916 739 17930 791
rect 17710 730 17930 739
rect 17850 720 17930 730
rect 17710 661 17790 680
rect 17710 609 17724 661
rect 17776 660 17790 661
rect 17776 610 17930 660
rect 17776 609 17790 610
rect 17710 590 17790 609
rect 17850 531 17930 550
rect 17850 530 17864 531
rect 17710 480 17864 530
rect 17850 479 17864 480
rect 17916 479 17930 531
rect 17850 460 17930 479
rect 17710 401 17790 420
rect 17710 349 17724 401
rect 17776 400 17790 401
rect 17960 400 18020 4310
rect 18270 4310 18670 4370
rect 18270 400 18330 4310
rect 18500 4241 18580 4260
rect 18500 4240 18514 4241
rect 18360 4234 18514 4240
rect 18360 4200 18430 4234
rect 18500 4200 18514 4234
rect 18360 4194 18514 4200
rect 18360 4190 18430 4194
rect 18500 4189 18514 4194
rect 18566 4189 18580 4241
rect 18500 4170 18580 4189
rect 18360 4112 18440 4130
rect 18360 4111 18571 4112
rect 18360 4059 18374 4111
rect 18426 4110 18571 4111
rect 18426 4060 18580 4110
rect 18426 4059 18440 4060
rect 18360 4040 18440 4059
rect 18500 3990 18580 4000
rect 18360 3981 18580 3990
rect 18360 3940 18514 3981
rect 18371 3938 18514 3940
rect 18500 3929 18514 3938
rect 18566 3929 18580 3981
rect 18500 3910 18580 3929
rect 18360 3861 18440 3880
rect 18360 3809 18374 3861
rect 18426 3860 18440 3861
rect 18426 3810 18580 3860
rect 18426 3809 18440 3810
rect 18360 3790 18440 3809
rect 18500 3731 18580 3750
rect 18500 3730 18514 3731
rect 18360 3680 18514 3730
rect 18500 3679 18514 3680
rect 18566 3679 18580 3731
rect 18500 3660 18580 3679
rect 18360 3601 18440 3620
rect 18360 3549 18374 3601
rect 18426 3600 18440 3601
rect 18426 3550 18580 3600
rect 18426 3549 18440 3550
rect 18360 3530 18440 3549
rect 18500 3472 18580 3490
rect 18371 3471 18580 3472
rect 18371 3470 18514 3471
rect 18360 3420 18514 3470
rect 18500 3419 18514 3420
rect 18566 3419 18580 3471
rect 18500 3400 18580 3419
rect 18360 3351 18440 3370
rect 18360 3299 18374 3351
rect 18426 3350 18440 3351
rect 18426 3300 18580 3350
rect 18426 3299 18571 3300
rect 18360 3298 18571 3299
rect 18360 3280 18440 3298
rect 18500 3221 18580 3240
rect 18500 3220 18514 3221
rect 18360 3170 18514 3220
rect 18500 3169 18514 3170
rect 18566 3169 18580 3221
rect 18500 3150 18580 3169
rect 18360 3091 18440 3110
rect 18360 3039 18374 3091
rect 18426 3090 18440 3091
rect 18426 3040 18580 3090
rect 18426 3039 18440 3040
rect 18360 3020 18440 3039
rect 18500 2961 18580 2980
rect 18500 2960 18514 2961
rect 18360 2910 18514 2960
rect 18500 2909 18514 2910
rect 18566 2909 18580 2961
rect 18500 2890 18580 2909
rect 18360 2832 18440 2850
rect 18360 2831 18571 2832
rect 18360 2779 18374 2831
rect 18426 2830 18571 2831
rect 18426 2780 18580 2830
rect 18426 2779 18440 2780
rect 18360 2760 18440 2779
rect 18500 2711 18580 2730
rect 18500 2710 18514 2711
rect 18360 2659 18514 2710
rect 18566 2659 18580 2711
rect 18360 2650 18580 2659
rect 18500 2640 18580 2650
rect 18360 2581 18440 2600
rect 18360 2529 18374 2581
rect 18426 2580 18440 2581
rect 18426 2530 18580 2580
rect 18426 2529 18440 2530
rect 18360 2510 18440 2529
rect 18500 2451 18580 2470
rect 18500 2450 18514 2451
rect 18360 2400 18514 2450
rect 18500 2399 18514 2400
rect 18566 2399 18580 2451
rect 18500 2380 18580 2399
rect 18360 2321 18440 2340
rect 18360 2269 18374 2321
rect 18426 2320 18440 2321
rect 18426 2270 18580 2320
rect 18426 2269 18440 2270
rect 18360 2250 18440 2269
rect 18500 2200 18580 2210
rect 18360 2191 18580 2200
rect 18360 2140 18514 2191
rect 18500 2139 18514 2140
rect 18566 2139 18580 2191
rect 18500 2120 18580 2139
rect 18360 2071 18440 2090
rect 18360 2019 18374 2071
rect 18426 2070 18440 2071
rect 18426 2019 18580 2070
rect 18360 2010 18580 2019
rect 18360 2000 18440 2010
rect 18500 1941 18580 1960
rect 18500 1940 18514 1941
rect 18360 1890 18514 1940
rect 18500 1889 18514 1890
rect 18566 1889 18580 1941
rect 18500 1870 18580 1889
rect 18360 1811 18440 1830
rect 18360 1759 18374 1811
rect 18426 1810 18440 1811
rect 18426 1760 18580 1810
rect 18426 1759 18440 1760
rect 18360 1740 18440 1759
rect 18500 1681 18580 1700
rect 18500 1680 18514 1681
rect 18360 1630 18514 1680
rect 18500 1629 18514 1630
rect 18566 1629 18580 1681
rect 18500 1610 18580 1629
rect 18360 1552 18440 1570
rect 18360 1551 18571 1552
rect 18360 1499 18374 1551
rect 18426 1550 18571 1551
rect 18426 1510 18580 1550
rect 18426 1506 18571 1510
rect 18426 1499 18440 1506
rect 18360 1480 18440 1499
rect 18500 1430 18580 1440
rect 18360 1421 18580 1430
rect 18360 1380 18514 1421
rect 18371 1378 18514 1380
rect 18500 1369 18514 1378
rect 18566 1369 18580 1421
rect 18500 1350 18580 1369
rect 18360 1301 18440 1320
rect 18360 1249 18374 1301
rect 18426 1300 18440 1301
rect 18610 1310 18670 4310
rect 19200 2213 19770 4790
rect 19200 1841 19262 2213
rect 19698 1841 19770 2213
rect 20070 1845 20130 6160
rect 20160 6116 20250 6130
rect 20160 6064 20179 6116
rect 20231 6110 20250 6116
rect 20231 6070 20380 6110
rect 20231 6064 20250 6070
rect 20160 6050 20250 6064
rect 20290 5986 20380 6000
rect 20290 5980 20309 5986
rect 20160 5940 20309 5980
rect 20290 5934 20309 5940
rect 20361 5934 20380 5986
rect 20290 5920 20380 5934
rect 20160 5856 20250 5870
rect 20160 5804 20179 5856
rect 20231 5850 20250 5856
rect 20231 5810 20380 5850
rect 20231 5804 20250 5810
rect 20160 5790 20250 5804
rect 20290 5726 20380 5740
rect 20290 5720 20309 5726
rect 20160 5680 20309 5720
rect 20290 5674 20309 5680
rect 20361 5674 20380 5726
rect 20290 5660 20380 5674
rect 20160 5606 20250 5620
rect 20160 5554 20179 5606
rect 20231 5600 20250 5606
rect 20231 5554 20380 5600
rect 20160 5550 20380 5554
rect 20160 5540 20250 5550
rect 20290 5476 20380 5490
rect 20290 5470 20309 5476
rect 20160 5424 20309 5470
rect 20361 5424 20380 5476
rect 20160 5420 20380 5424
rect 20290 5410 20380 5420
rect 20160 5346 20250 5360
rect 20160 5294 20179 5346
rect 20231 5340 20250 5346
rect 20231 5300 20380 5340
rect 20231 5294 20250 5300
rect 20160 5280 20250 5294
rect 20290 5216 20380 5230
rect 20290 5210 20309 5216
rect 20160 5170 20309 5210
rect 20290 5164 20309 5170
rect 20361 5164 20380 5216
rect 20290 5150 20380 5164
rect 20160 5090 20250 5100
rect 20160 5086 20380 5090
rect 20160 5034 20179 5086
rect 20231 5040 20380 5086
rect 20231 5034 20250 5040
rect 20160 5020 20250 5034
rect 20290 4960 20380 4970
rect 20160 4956 20380 4960
rect 20160 4910 20309 4956
rect 20290 4904 20309 4910
rect 20361 4904 20380 4956
rect 20290 4890 20380 4904
rect 20160 4830 20250 4840
rect 20160 4826 20380 4830
rect 20160 4774 20179 4826
rect 20231 4780 20380 4826
rect 20231 4774 20250 4780
rect 20160 4760 20250 4774
rect 20290 4706 20380 4720
rect 20290 4700 20309 4706
rect 20160 4660 20309 4700
rect 20290 4654 20309 4660
rect 20361 4654 20380 4706
rect 20290 4640 20380 4654
rect 20160 4576 20250 4590
rect 20160 4524 20179 4576
rect 20231 4570 20250 4576
rect 20231 4530 20380 4570
rect 20231 4524 20250 4530
rect 20160 4510 20250 4524
rect 20290 4446 20380 4460
rect 20290 4440 20309 4446
rect 20160 4400 20309 4440
rect 20290 4394 20309 4400
rect 20361 4394 20380 4446
rect 20290 4380 20380 4394
rect 20160 4320 20250 4330
rect 20160 4316 20380 4320
rect 20160 4264 20179 4316
rect 20231 4270 20380 4316
rect 20231 4264 20250 4270
rect 20160 4250 20250 4264
rect 20290 4196 20380 4210
rect 20290 4190 20309 4196
rect 20160 4144 20309 4190
rect 20361 4144 20380 4196
rect 20160 4140 20380 4144
rect 20290 4130 20380 4140
rect 20290 3865 20380 3875
rect 20160 3861 20380 3865
rect 20160 3815 20309 3861
rect 20290 3809 20309 3815
rect 20361 3809 20380 3861
rect 20290 3795 20380 3809
rect 20160 3741 20250 3755
rect 20160 3689 20179 3741
rect 20231 3735 20250 3741
rect 20231 3689 20380 3735
rect 20160 3685 20380 3689
rect 20160 3675 20250 3685
rect 20290 3611 20380 3625
rect 20290 3605 20309 3611
rect 20160 3565 20309 3605
rect 20169 3559 20309 3565
rect 20361 3559 20380 3611
rect 20290 3545 20380 3559
rect 20160 3481 20250 3495
rect 20160 3429 20179 3481
rect 20231 3477 20250 3481
rect 20231 3475 20369 3477
rect 20231 3435 20380 3475
rect 20231 3431 20369 3435
rect 20231 3429 20250 3431
rect 20160 3415 20250 3429
rect 20290 3351 20380 3365
rect 20290 3349 20309 3351
rect 20169 3345 20309 3349
rect 20160 3305 20309 3345
rect 20169 3303 20309 3305
rect 20290 3299 20309 3303
rect 20361 3299 20380 3351
rect 20290 3285 20380 3299
rect 20160 3231 20250 3245
rect 20160 3179 20179 3231
rect 20231 3225 20250 3231
rect 20231 3179 20380 3225
rect 20160 3175 20380 3179
rect 20160 3165 20250 3175
rect 20290 3101 20380 3115
rect 20290 3095 20309 3101
rect 20160 3049 20309 3095
rect 20361 3049 20380 3101
rect 20160 3045 20380 3049
rect 20290 3035 20380 3045
rect 20160 2971 20250 2985
rect 20160 2919 20179 2971
rect 20231 2965 20250 2971
rect 20231 2919 20380 2965
rect 20160 2915 20380 2919
rect 20160 2905 20250 2915
rect 20290 2841 20380 2855
rect 20290 2837 20309 2841
rect 20169 2835 20309 2837
rect 20160 2795 20309 2835
rect 20169 2791 20309 2795
rect 20290 2789 20309 2791
rect 20361 2789 20380 2841
rect 20290 2775 20380 2789
rect 20160 2711 20250 2725
rect 20160 2659 20179 2711
rect 20231 2709 20250 2711
rect 20231 2705 20369 2709
rect 20231 2665 20380 2705
rect 20231 2663 20369 2665
rect 20231 2659 20250 2663
rect 20160 2645 20250 2659
rect 20290 2585 20380 2595
rect 20160 2581 20380 2585
rect 20160 2535 20309 2581
rect 20290 2529 20309 2535
rect 20361 2529 20380 2581
rect 20290 2515 20380 2529
rect 20160 2455 20250 2465
rect 20160 2451 20380 2455
rect 20160 2399 20179 2451
rect 20231 2405 20380 2451
rect 20231 2399 20250 2405
rect 20160 2385 20250 2399
rect 20290 2331 20380 2345
rect 20290 2325 20309 2331
rect 20160 2285 20309 2325
rect 20169 2279 20309 2285
rect 20361 2279 20380 2331
rect 20290 2265 20380 2279
rect 20160 2201 20250 2215
rect 20160 2149 20179 2201
rect 20231 2197 20250 2201
rect 20231 2195 20369 2197
rect 20231 2155 20380 2195
rect 20231 2151 20369 2155
rect 20231 2149 20250 2151
rect 20160 2135 20250 2149
rect 20290 2071 20380 2085
rect 20290 2069 20309 2071
rect 20169 2065 20309 2069
rect 20160 2025 20309 2065
rect 20169 2023 20309 2025
rect 20290 2019 20309 2023
rect 20361 2019 20380 2071
rect 20290 2005 20380 2019
rect 20160 1941 20250 1955
rect 20160 1889 20179 1941
rect 20231 1935 20369 1941
rect 20231 1895 20380 1935
rect 20231 1889 20250 1895
rect 20160 1875 20250 1889
rect 20410 1845 20470 6160
rect 20820 5520 21340 5580
rect 20820 4180 20880 5520
rect 20910 5476 21000 5490
rect 20910 5424 20929 5476
rect 20981 5470 21000 5476
rect 20981 5424 21130 5470
rect 20910 5420 21130 5424
rect 20910 5410 21000 5420
rect 21040 5346 21130 5360
rect 21040 5340 21059 5346
rect 20910 5294 21059 5340
rect 21111 5294 21130 5346
rect 20910 5290 21130 5294
rect 21040 5280 21130 5290
rect 20910 5220 21000 5230
rect 20910 5216 21130 5220
rect 20910 5164 20929 5216
rect 20981 5170 21130 5216
rect 20981 5164 21000 5170
rect 20910 5150 21000 5164
rect 21040 5091 21130 5110
rect 21040 5090 21059 5091
rect 20910 5040 21059 5090
rect 21040 5039 21059 5040
rect 21111 5039 21130 5091
rect 21040 5020 21130 5039
rect 20910 4966 21000 4980
rect 20910 4914 20929 4966
rect 20981 4960 21000 4966
rect 20981 4914 21130 4960
rect 20910 4910 21130 4914
rect 20910 4900 21000 4910
rect 21040 4836 21130 4850
rect 21040 4830 21059 4836
rect 20910 4784 21059 4830
rect 21111 4784 21130 4836
rect 20910 4780 21130 4784
rect 21040 4770 21130 4780
rect 20910 4706 21000 4720
rect 20910 4654 20929 4706
rect 20981 4700 21000 4706
rect 20981 4660 21130 4700
rect 20981 4654 21000 4660
rect 20910 4640 21000 4654
rect 21040 4576 21130 4590
rect 21040 4570 21059 4576
rect 20910 4530 21059 4570
rect 21040 4524 21059 4530
rect 21111 4524 21130 4576
rect 21040 4510 21130 4524
rect 20910 4450 21000 4460
rect 20910 4446 21130 4450
rect 20910 4394 20929 4446
rect 20981 4400 21130 4446
rect 20981 4394 21000 4400
rect 20910 4380 21000 4394
rect 21040 4320 21130 4330
rect 20910 4316 21130 4320
rect 20910 4270 21059 4316
rect 21040 4264 21059 4270
rect 21111 4264 21130 4316
rect 21040 4250 21130 4264
rect 20910 4196 21000 4210
rect 20910 4144 20929 4196
rect 20981 4190 21000 4196
rect 20981 4144 21130 4190
rect 21160 4180 21220 5520
rect 20910 4140 21130 4144
rect 20910 4130 21000 4140
rect 20910 3875 21000 3885
rect 20910 3871 21130 3875
rect 20820 2495 20880 3835
rect 20910 3819 20929 3871
rect 20981 3825 21130 3871
rect 20981 3819 21000 3825
rect 20910 3805 21000 3819
rect 21040 3751 21130 3765
rect 21040 3745 21059 3751
rect 20910 3699 21059 3745
rect 21111 3699 21130 3751
rect 20910 3695 21130 3699
rect 21040 3685 21130 3695
rect 20910 3621 21000 3635
rect 20910 3569 20929 3621
rect 20981 3615 21000 3621
rect 20981 3569 21130 3615
rect 20910 3565 21130 3569
rect 20910 3555 21000 3565
rect 21040 3491 21130 3505
rect 21040 3487 21059 3491
rect 20919 3485 21059 3487
rect 20910 3445 21059 3485
rect 20919 3441 21059 3445
rect 21040 3439 21059 3441
rect 21111 3439 21130 3491
rect 21040 3425 21130 3439
rect 20910 3361 21000 3375
rect 20910 3309 20929 3361
rect 20981 3359 21000 3361
rect 20981 3355 21119 3359
rect 20981 3315 21130 3355
rect 20981 3313 21119 3315
rect 20981 3309 21000 3313
rect 20910 3295 21000 3309
rect 21040 3235 21130 3245
rect 20910 3231 21130 3235
rect 20910 3185 21059 3231
rect 21040 3179 21059 3185
rect 21111 3179 21130 3231
rect 21040 3165 21130 3179
rect 20910 3105 21000 3115
rect 20910 3101 21130 3105
rect 20910 3049 20929 3101
rect 20981 3055 21130 3101
rect 20981 3049 21000 3055
rect 20910 3035 21000 3049
rect 21040 2976 21130 2995
rect 21040 2975 21059 2976
rect 20910 2925 21059 2975
rect 21040 2924 21059 2925
rect 21111 2924 21130 2976
rect 21040 2905 21130 2924
rect 20910 2851 21000 2865
rect 20910 2799 20929 2851
rect 20981 2847 21000 2851
rect 20981 2845 21119 2847
rect 20981 2799 21130 2845
rect 20910 2795 21130 2799
rect 20910 2785 21000 2795
rect 21040 2725 21130 2735
rect 20910 2721 21130 2725
rect 20910 2675 21059 2721
rect 20919 2673 21059 2675
rect 21040 2669 21059 2673
rect 21111 2669 21130 2721
rect 21040 2655 21130 2669
rect 20910 2595 21000 2605
rect 20910 2591 21130 2595
rect 20910 2539 20929 2591
rect 20981 2545 21130 2591
rect 20981 2539 21000 2545
rect 20910 2525 21000 2539
rect 21160 2495 21220 3835
rect 20820 2435 21340 2495
rect 19200 1800 19770 1841
rect 18426 1250 18580 1300
rect 18610 1280 19240 1310
rect 18426 1249 18440 1250
rect 18360 1230 18440 1249
rect 18610 1249 19750 1280
rect 18500 1171 18580 1190
rect 18500 1170 18514 1171
rect 18360 1120 18514 1170
rect 18500 1119 18514 1120
rect 18566 1119 18580 1171
rect 18500 1100 18580 1119
rect 18360 1041 18440 1060
rect 18360 989 18374 1041
rect 18426 1040 18440 1041
rect 18426 990 18580 1040
rect 18426 989 18440 990
rect 18360 970 18440 989
rect 18610 941 19245 1249
rect 19745 941 19750 1249
rect 18500 912 18580 930
rect 18371 911 18580 912
rect 18371 910 18514 911
rect 18360 860 18514 910
rect 18500 859 18514 860
rect 18566 859 18580 911
rect 18500 840 18580 859
rect 18610 910 19750 941
rect 18610 880 19240 910
rect 18360 791 18440 810
rect 18360 739 18374 791
rect 18426 790 18440 791
rect 18426 739 18580 790
rect 18360 730 18580 739
rect 18360 720 18440 730
rect 18500 661 18580 680
rect 18500 660 18514 661
rect 18360 610 18514 660
rect 18500 609 18514 610
rect 18566 609 18580 661
rect 18500 590 18580 609
rect 18360 531 18440 550
rect 18360 479 18374 531
rect 18426 530 18440 531
rect 18426 480 18580 530
rect 18426 479 18440 480
rect 18360 460 18440 479
rect 18500 401 18580 420
rect 18500 400 18514 401
rect 17776 350 17930 400
rect 18360 350 18514 400
rect 17776 349 17790 350
rect 17710 330 17790 349
rect 18500 349 18514 350
rect 18566 349 18580 401
rect 18610 400 18670 880
rect 18500 330 18580 349
rect 17390 -132 17495 -125
rect 17390 -160 17414 -132
rect 16985 -184 17414 -160
rect 17466 -160 17495 -132
rect 17775 -137 17880 -120
rect 17775 -160 17799 -137
rect 17466 -184 17799 -160
rect 16985 -189 17799 -184
rect 17851 -160 17880 -137
rect 17980 -132 18085 -120
rect 17980 -160 18009 -132
rect 17851 -184 18009 -160
rect 18061 -160 18085 -132
rect 18061 -184 19305 -160
rect 17851 -189 19305 -184
rect 16985 -210 19305 -189
rect 16985 -365 17040 -240
rect 17070 -252 17145 -240
rect 17070 -304 17081 -252
rect 17133 -304 17145 -252
rect 17070 -315 17145 -304
rect 16970 -377 17045 -365
rect 16970 -429 16981 -377
rect 17033 -429 17045 -377
rect 16970 -440 17045 -429
rect 17080 -440 17135 -315
rect 17175 -365 17230 -240
rect 17260 -252 17335 -240
rect 17260 -304 17271 -252
rect 17323 -304 17335 -252
rect 17260 -315 17335 -304
rect 17165 -377 17240 -365
rect 17165 -429 17176 -377
rect 17228 -429 17240 -377
rect 17165 -440 17240 -429
rect 17275 -440 17325 -315
rect 17370 -365 17425 -240
rect 17455 -252 17530 -240
rect 17455 -304 17466 -252
rect 17518 -304 17530 -252
rect 17455 -315 17530 -304
rect 17360 -377 17435 -365
rect 17360 -429 17371 -377
rect 17423 -429 17435 -377
rect 17360 -440 17435 -429
rect 17465 -440 17520 -315
rect 17560 -365 17615 -240
rect 17645 -252 17720 -240
rect 17645 -304 17656 -252
rect 17708 -304 17720 -252
rect 17645 -315 17720 -304
rect 17550 -377 17625 -365
rect 17550 -429 17561 -377
rect 17613 -429 17625 -377
rect 17550 -440 17625 -429
rect 17655 -440 17710 -315
rect 17755 -365 17810 -240
rect 17840 -252 17915 -240
rect 17840 -304 17851 -252
rect 17903 -304 17915 -252
rect 17840 -315 17915 -304
rect 17740 -377 17815 -365
rect 17740 -429 17751 -377
rect 17803 -429 17815 -377
rect 17740 -440 17815 -429
rect 17850 -440 17905 -315
rect 17945 -365 18000 -240
rect 17935 -377 18010 -365
rect 17935 -429 17946 -377
rect 17998 -429 18010 -377
rect 17935 -440 18010 -429
rect 18125 -470 18165 -210
rect 18290 -365 18345 -240
rect 18375 -252 18450 -240
rect 18375 -304 18386 -252
rect 18438 -304 18450 -252
rect 18375 -315 18450 -304
rect 18280 -377 18355 -365
rect 18280 -429 18291 -377
rect 18343 -429 18355 -377
rect 18280 -440 18355 -429
rect 18385 -440 18440 -315
rect 18480 -365 18535 -240
rect 18570 -252 18645 -240
rect 18570 -304 18581 -252
rect 18633 -304 18645 -252
rect 18570 -315 18645 -304
rect 18475 -377 18550 -365
rect 18475 -429 18486 -377
rect 18538 -429 18550 -377
rect 18475 -440 18550 -429
rect 18580 -440 18635 -315
rect 18675 -365 18730 -240
rect 18760 -252 18835 -240
rect 18760 -304 18771 -252
rect 18823 -304 18835 -252
rect 18760 -315 18835 -304
rect 18665 -377 18740 -365
rect 18665 -429 18676 -377
rect 18728 -429 18740 -377
rect 18665 -440 18740 -429
rect 18770 -440 18825 -315
rect 18865 -365 18920 -240
rect 18955 -252 19030 -240
rect 18955 -304 18966 -252
rect 19018 -304 19030 -252
rect 18955 -315 19030 -304
rect 18855 -377 18930 -365
rect 18855 -429 18866 -377
rect 18918 -429 18930 -377
rect 18855 -440 18930 -429
rect 18965 -440 19015 -315
rect 19060 -365 19115 -240
rect 19145 -252 19220 -240
rect 19145 -304 19156 -252
rect 19208 -304 19220 -252
rect 19145 -315 19220 -304
rect 19050 -377 19125 -365
rect 19050 -429 19061 -377
rect 19113 -429 19125 -377
rect 19050 -440 19125 -429
rect 19155 -440 19210 -315
rect 19250 -365 19305 -240
rect 19245 -377 19320 -365
rect 19245 -429 19256 -377
rect 19308 -429 19320 -377
rect 19245 -440 19320 -429
rect 16980 -520 19310 -470
<< via1 >>
rect 17329 7054 17381 7106
rect 17459 6924 17511 6976
rect 17329 6794 17381 6846
rect 17459 6664 17511 6716
rect 17329 6534 17381 6586
rect 17459 6404 17511 6456
rect 17329 6274 17381 6326
rect 17459 6154 17511 6206
rect 17329 6024 17381 6076
rect 17459 5904 17511 5956
rect 17329 5774 17381 5826
rect 17459 5644 17511 5696
rect 17329 5514 17381 5566
rect 17459 5384 17511 5436
rect 17329 5254 17381 5306
rect 17979 7054 18031 7106
rect 18109 6924 18161 6976
rect 17979 6794 18031 6846
rect 18109 6664 18161 6716
rect 17979 6534 18031 6586
rect 18109 6404 18161 6456
rect 17979 6274 18031 6326
rect 18109 6154 18161 6206
rect 17979 6024 18031 6076
rect 18109 5904 18161 5956
rect 17979 5774 18031 5826
rect 18109 5644 18161 5696
rect 17979 5514 18031 5566
rect 18109 5384 18161 5436
rect 17979 5254 18031 5306
rect 18629 7054 18681 7106
rect 18759 6924 18811 6976
rect 18629 6794 18681 6846
rect 18759 6664 18811 6716
rect 18629 6534 18681 6586
rect 18759 6404 18811 6456
rect 18629 6274 18681 6326
rect 18759 6154 18811 6206
rect 18629 6024 18681 6076
rect 18759 5904 18811 5956
rect 18629 5774 18681 5826
rect 18759 5644 18811 5696
rect 18629 5514 18681 5566
rect 18759 5384 18811 5436
rect 18629 5254 18681 5306
rect 19237 6331 19737 6703
rect 17459 5124 17511 5176
rect 18109 5124 18161 5176
rect 18759 5124 18811 5176
rect 17724 4189 17776 4241
rect 17864 4059 17916 4111
rect 17724 3929 17776 3981
rect 17864 3809 17916 3861
rect 17724 3679 17776 3731
rect 17864 3549 17916 3601
rect 17724 3419 17776 3471
rect 17864 3299 17916 3351
rect 17724 3169 17776 3221
rect 17864 3039 17916 3091
rect 17724 2909 17776 2961
rect 17864 2779 17916 2831
rect 17724 2659 17776 2711
rect 17864 2529 17916 2581
rect 17724 2399 17776 2451
rect 17864 2269 17916 2321
rect 17724 2139 17776 2191
rect 17864 2019 17916 2071
rect 17724 1889 17776 1941
rect 17864 1759 17916 1811
rect 17724 1629 17776 1681
rect 17864 1499 17916 1551
rect 17724 1369 17776 1421
rect 17864 1249 17916 1301
rect 17724 1119 17776 1171
rect 17864 989 17916 1041
rect 17724 859 17776 911
rect 17864 739 17916 791
rect 17724 609 17776 661
rect 17864 479 17916 531
rect 17724 349 17776 401
rect 18514 4189 18566 4241
rect 18374 4059 18426 4111
rect 18514 3929 18566 3981
rect 18374 3809 18426 3861
rect 18514 3679 18566 3731
rect 18374 3549 18426 3601
rect 18514 3419 18566 3471
rect 18374 3299 18426 3351
rect 18514 3169 18566 3221
rect 18374 3039 18426 3091
rect 18514 2909 18566 2961
rect 18374 2779 18426 2831
rect 18514 2659 18566 2711
rect 18374 2529 18426 2581
rect 18514 2399 18566 2451
rect 18374 2269 18426 2321
rect 18514 2139 18566 2191
rect 18374 2019 18426 2071
rect 18514 1889 18566 1941
rect 18374 1759 18426 1811
rect 18514 1629 18566 1681
rect 18374 1499 18426 1551
rect 18514 1369 18566 1421
rect 18374 1249 18426 1301
rect 19262 1841 19698 2213
rect 20179 6064 20231 6116
rect 20309 5934 20361 5986
rect 20179 5804 20231 5856
rect 20309 5674 20361 5726
rect 20179 5554 20231 5606
rect 20309 5424 20361 5476
rect 20179 5294 20231 5346
rect 20309 5164 20361 5216
rect 20179 5034 20231 5086
rect 20309 4904 20361 4956
rect 20179 4774 20231 4826
rect 20309 4654 20361 4706
rect 20179 4524 20231 4576
rect 20309 4394 20361 4446
rect 20179 4264 20231 4316
rect 20309 4144 20361 4196
rect 20309 3809 20361 3861
rect 20179 3689 20231 3741
rect 20309 3559 20361 3611
rect 20179 3429 20231 3481
rect 20309 3299 20361 3351
rect 20179 3179 20231 3231
rect 20309 3049 20361 3101
rect 20179 2919 20231 2971
rect 20309 2789 20361 2841
rect 20179 2659 20231 2711
rect 20309 2529 20361 2581
rect 20179 2399 20231 2451
rect 20309 2279 20361 2331
rect 20179 2149 20231 2201
rect 20309 2019 20361 2071
rect 20179 1889 20231 1941
rect 20929 5424 20981 5476
rect 21059 5294 21111 5346
rect 20929 5164 20981 5216
rect 21059 5039 21111 5091
rect 20929 4914 20981 4966
rect 21059 4784 21111 4836
rect 20929 4654 20981 4706
rect 21059 4524 21111 4576
rect 20929 4394 20981 4446
rect 21059 4264 21111 4316
rect 20929 4144 20981 4196
rect 20929 3819 20981 3871
rect 21059 3699 21111 3751
rect 20929 3569 20981 3621
rect 21059 3439 21111 3491
rect 20929 3309 20981 3361
rect 21059 3179 21111 3231
rect 20929 3049 20981 3101
rect 21059 2924 21111 2976
rect 20929 2799 20981 2851
rect 21059 2669 21111 2721
rect 20929 2539 20981 2591
rect 18514 1119 18566 1171
rect 18374 989 18426 1041
rect 19245 941 19745 1249
rect 18514 859 18566 911
rect 18374 739 18426 791
rect 18514 609 18566 661
rect 18374 479 18426 531
rect 18514 349 18566 401
rect 17414 -184 17466 -132
rect 17799 -189 17851 -137
rect 18009 -184 18061 -132
rect 17081 -304 17133 -252
rect 16981 -429 17033 -377
rect 17271 -304 17323 -252
rect 17176 -429 17228 -377
rect 17466 -304 17518 -252
rect 17371 -429 17423 -377
rect 17656 -304 17708 -252
rect 17561 -429 17613 -377
rect 17851 -304 17903 -252
rect 17751 -429 17803 -377
rect 17946 -429 17998 -377
rect 18386 -304 18438 -252
rect 18291 -429 18343 -377
rect 18581 -304 18633 -252
rect 18486 -429 18538 -377
rect 18771 -304 18823 -252
rect 18676 -429 18728 -377
rect 18966 -304 19018 -252
rect 18866 -429 18918 -377
rect 19156 -304 19208 -252
rect 19061 -429 19113 -377
rect 19256 -429 19308 -377
<< metal2 >>
rect 17440 7235 17720 7275
rect 17440 7179 17469 7235
rect 17525 7179 17549 7235
rect 17605 7179 17629 7235
rect 17685 7179 17720 7235
rect 17100 7106 17400 7120
rect 17100 7054 17329 7106
rect 17381 7054 17400 7106
rect 17100 6846 17400 7054
rect 17100 6794 17329 6846
rect 17381 6794 17400 6846
rect 17100 6586 17400 6794
rect 17100 6534 17329 6586
rect 17381 6534 17400 6586
rect 17100 6326 17400 6534
rect 17100 6274 17329 6326
rect 17381 6274 17400 6326
rect 17100 6076 17400 6274
rect 17100 6024 17329 6076
rect 17381 6024 17400 6076
rect 17100 5826 17400 6024
rect 17100 5774 17329 5826
rect 17381 5774 17400 5826
rect 17100 5566 17400 5774
rect 17100 5514 17329 5566
rect 17381 5514 17400 5566
rect 17100 5306 17400 5514
rect 17100 5254 17329 5306
rect 17381 5254 17400 5306
rect 17100 5000 17400 5254
rect 17440 6976 17720 7179
rect 18090 7235 18370 7275
rect 18090 7179 18124 7235
rect 18180 7179 18204 7235
rect 18260 7179 18284 7235
rect 18340 7179 18370 7235
rect 17440 6924 17459 6976
rect 17511 6924 17720 6976
rect 17440 6716 17720 6924
rect 17440 6664 17459 6716
rect 17511 6664 17720 6716
rect 17440 6456 17720 6664
rect 17440 6404 17459 6456
rect 17511 6404 17720 6456
rect 17440 6206 17720 6404
rect 17440 6154 17459 6206
rect 17511 6154 17720 6206
rect 17440 5956 17720 6154
rect 17440 5904 17459 5956
rect 17511 5904 17720 5956
rect 17440 5696 17720 5904
rect 17440 5644 17459 5696
rect 17511 5644 17720 5696
rect 17440 5436 17720 5644
rect 17440 5384 17459 5436
rect 17511 5384 17720 5436
rect 17440 5176 17720 5384
rect 17440 5124 17459 5176
rect 17511 5124 17720 5176
rect 17440 5110 17720 5124
rect 17760 7106 18050 7120
rect 17760 7054 17979 7106
rect 18031 7054 18050 7106
rect 17760 6846 18050 7054
rect 17760 6794 17979 6846
rect 18031 6794 18050 6846
rect 17760 6586 18050 6794
rect 17760 6534 17979 6586
rect 18031 6534 18050 6586
rect 17760 6326 18050 6534
rect 17760 6274 17979 6326
rect 18031 6274 18050 6326
rect 17760 6076 18050 6274
rect 17760 6024 17979 6076
rect 18031 6024 18050 6076
rect 17760 5826 18050 6024
rect 17760 5774 17979 5826
rect 18031 5774 18050 5826
rect 17760 5566 18050 5774
rect 17760 5514 17979 5566
rect 18031 5514 18050 5566
rect 17760 5306 18050 5514
rect 17760 5254 17979 5306
rect 18031 5254 18050 5306
rect 17760 5000 18050 5254
rect 18090 6976 18370 7179
rect 18740 7235 19020 7275
rect 18740 7179 18769 7235
rect 18825 7179 18849 7235
rect 18905 7179 18929 7235
rect 18985 7179 19020 7235
rect 18090 6924 18109 6976
rect 18161 6924 18370 6976
rect 18090 6716 18370 6924
rect 18090 6664 18109 6716
rect 18161 6664 18370 6716
rect 18090 6456 18370 6664
rect 18090 6404 18109 6456
rect 18161 6404 18370 6456
rect 18090 6206 18370 6404
rect 18090 6154 18109 6206
rect 18161 6154 18370 6206
rect 18090 5956 18370 6154
rect 18090 5904 18109 5956
rect 18161 5904 18370 5956
rect 18090 5696 18370 5904
rect 18090 5644 18109 5696
rect 18161 5644 18370 5696
rect 18090 5436 18370 5644
rect 18090 5384 18109 5436
rect 18161 5384 18370 5436
rect 18090 5176 18370 5384
rect 18090 5124 18109 5176
rect 18161 5124 18370 5176
rect 18090 5110 18370 5124
rect 18410 7106 18700 7120
rect 18410 7054 18629 7106
rect 18681 7054 18700 7106
rect 18410 6846 18700 7054
rect 18410 6794 18629 6846
rect 18681 6794 18700 6846
rect 18410 6586 18700 6794
rect 18410 6534 18629 6586
rect 18681 6534 18700 6586
rect 18410 6326 18700 6534
rect 18410 6274 18629 6326
rect 18681 6274 18700 6326
rect 18410 6076 18700 6274
rect 18410 6024 18629 6076
rect 18681 6024 18700 6076
rect 18410 5826 18700 6024
rect 18410 5774 18629 5826
rect 18681 5774 18700 5826
rect 18410 5566 18700 5774
rect 18410 5514 18629 5566
rect 18681 5514 18700 5566
rect 18410 5306 18700 5514
rect 18410 5254 18629 5306
rect 18681 5254 18700 5306
rect 18410 5000 18700 5254
rect 18740 6976 19020 7179
rect 18740 6924 18759 6976
rect 18811 6924 19020 6976
rect 18740 6716 19020 6924
rect 18740 6664 18759 6716
rect 18811 6664 19020 6716
rect 18740 6456 19020 6664
rect 18740 6404 18759 6456
rect 18811 6404 19020 6456
rect 18740 6206 19020 6404
rect 19210 6703 21340 6745
rect 19210 6331 19237 6703
rect 19737 6331 21340 6703
rect 19210 6300 21340 6331
rect 18740 6154 18759 6206
rect 18811 6154 19020 6206
rect 18740 5956 19020 6154
rect 18740 5904 18759 5956
rect 18811 5904 19020 5956
rect 18740 5696 19020 5904
rect 18740 5644 18759 5696
rect 18811 5644 19020 5696
rect 18740 5436 19020 5644
rect 18740 5384 18759 5436
rect 18811 5384 19020 5436
rect 18740 5176 19020 5384
rect 18740 5124 18759 5176
rect 18811 5124 19020 5176
rect 18740 5110 19020 5124
rect 19950 6116 20250 6150
rect 19950 6098 20179 6116
rect 19950 5962 19992 6098
rect 20231 6064 20250 6116
rect 20208 5962 20250 6064
rect 19950 5856 20250 5962
rect 19950 5804 20179 5856
rect 20231 5804 20250 5856
rect 19950 5606 20250 5804
rect 19950 5554 20179 5606
rect 20231 5554 20250 5606
rect 19950 5346 20250 5554
rect 19950 5294 20179 5346
rect 20231 5294 20250 5346
rect 17100 4400 18700 5000
rect 19950 5086 20250 5294
rect 19950 5034 20179 5086
rect 20231 5034 20250 5086
rect 19950 4826 20250 5034
rect 19950 4774 20179 4826
rect 20231 4774 20250 4826
rect 19950 4576 20250 4774
rect 19950 4524 20179 4576
rect 20231 4524 20250 4576
rect 17190 4241 17790 4260
rect 17190 4189 17724 4241
rect 17776 4189 17790 4241
rect 17190 3981 17790 4189
rect 17190 3929 17724 3981
rect 17776 3929 17790 3981
rect 17190 3731 17790 3929
rect 17190 3679 17724 3731
rect 17776 3679 17790 3731
rect 17190 3471 17790 3679
rect 17190 3419 17724 3471
rect 17776 3419 17790 3471
rect 17190 3221 17790 3419
rect 17190 3169 17724 3221
rect 17776 3169 17790 3221
rect 17190 2961 17790 3169
rect 17190 2909 17724 2961
rect 17776 2909 17790 2961
rect 17190 2711 17790 2909
rect 17190 2659 17724 2711
rect 17776 2659 17790 2711
rect 17190 2451 17790 2659
rect 17190 2399 17724 2451
rect 17776 2399 17790 2451
rect 17190 2191 17790 2399
rect 17190 2139 17724 2191
rect 17776 2139 17790 2191
rect 17190 1941 17790 2139
rect 17190 1889 17724 1941
rect 17776 1889 17790 1941
rect 17190 1681 17790 1889
rect 17190 1629 17724 1681
rect 17776 1629 17790 1681
rect 17190 1421 17790 1629
rect 17190 1369 17724 1421
rect 17776 1369 17790 1421
rect 17190 1171 17790 1369
rect 17190 1119 17724 1171
rect 17776 1119 17790 1171
rect 17190 911 17790 1119
rect 17190 859 17724 911
rect 17776 859 17790 911
rect 17190 661 17790 859
rect 17190 609 17724 661
rect 17776 609 17790 661
rect 17190 401 17790 609
rect 17850 4111 18440 4400
rect 19950 4316 20250 4524
rect 19950 4264 20179 4316
rect 20231 4264 20250 4316
rect 17850 4059 17864 4111
rect 17916 4059 18374 4111
rect 18426 4059 18440 4111
rect 17850 3861 18440 4059
rect 17850 3809 17864 3861
rect 17916 3809 18374 3861
rect 18426 3809 18440 3861
rect 17850 3601 18440 3809
rect 17850 3549 17864 3601
rect 17916 3549 18374 3601
rect 18426 3549 18440 3601
rect 17850 3351 18440 3549
rect 17850 3299 17864 3351
rect 17916 3299 18374 3351
rect 18426 3299 18440 3351
rect 17850 3091 18440 3299
rect 17850 3039 17864 3091
rect 17916 3039 18374 3091
rect 18426 3039 18440 3091
rect 17850 2831 18440 3039
rect 17850 2779 17864 2831
rect 17916 2779 18374 2831
rect 18426 2779 18440 2831
rect 17850 2581 18440 2779
rect 17850 2529 17864 2581
rect 17916 2529 18374 2581
rect 18426 2529 18440 2581
rect 17850 2321 18440 2529
rect 17850 2269 17864 2321
rect 17916 2269 18374 2321
rect 18426 2269 18440 2321
rect 17850 2071 18440 2269
rect 17850 2019 17864 2071
rect 17916 2019 18374 2071
rect 18426 2019 18440 2071
rect 17850 1811 18440 2019
rect 17850 1759 17864 1811
rect 17916 1759 18374 1811
rect 18426 1759 18440 1811
rect 17850 1551 18440 1759
rect 17850 1499 17864 1551
rect 17916 1499 18374 1551
rect 18426 1499 18440 1551
rect 17850 1301 18440 1499
rect 17850 1249 17864 1301
rect 17916 1249 18374 1301
rect 18426 1249 18440 1301
rect 17850 1041 18440 1249
rect 17850 989 17864 1041
rect 17916 989 18374 1041
rect 18426 989 18440 1041
rect 17850 791 18440 989
rect 17850 739 17864 791
rect 17916 739 18374 791
rect 18426 739 18440 791
rect 17850 531 18440 739
rect 17850 479 17864 531
rect 17916 479 18374 531
rect 18426 479 18440 531
rect 17850 460 18440 479
rect 18500 4241 19100 4260
rect 18500 4189 18514 4241
rect 18566 4189 19100 4241
rect 18500 3981 19100 4189
rect 18500 3929 18514 3981
rect 18566 3929 19100 3981
rect 18500 3731 19100 3929
rect 18500 3679 18514 3731
rect 18566 3679 19100 3731
rect 18500 3471 19100 3679
rect 18500 3419 18514 3471
rect 18566 3419 19100 3471
rect 18500 3221 19100 3419
rect 18500 3169 18514 3221
rect 18566 3169 19100 3221
rect 18500 2961 19100 3169
rect 18500 2909 18514 2961
rect 18566 2909 19100 2961
rect 18500 2711 19100 2909
rect 18500 2659 18514 2711
rect 18566 2659 19100 2711
rect 18500 2451 19100 2659
rect 18500 2399 18514 2451
rect 18566 2399 19100 2451
rect 18500 2191 19100 2399
rect 19950 3741 20250 4264
rect 19950 3689 20179 3741
rect 20231 3689 20250 3741
rect 19950 3481 20250 3689
rect 19950 3429 20179 3481
rect 20231 3429 20250 3481
rect 19950 3231 20250 3429
rect 19950 3179 20179 3231
rect 20231 3179 20250 3231
rect 19950 2971 20250 3179
rect 19950 2919 20179 2971
rect 20231 2919 20250 2971
rect 19950 2711 20250 2919
rect 19950 2659 20179 2711
rect 20231 2659 20250 2711
rect 19950 2451 20250 2659
rect 19950 2399 20179 2451
rect 20231 2399 20250 2451
rect 18500 2139 18514 2191
rect 18566 2139 19100 2191
rect 18500 1941 19100 2139
rect 18500 1889 18514 1941
rect 18566 1889 19100 1941
rect 18500 1681 19100 1889
rect 19200 2213 19770 2255
rect 19200 2175 19262 2213
rect 19698 2175 19770 2213
rect 19200 1879 19252 2175
rect 19708 1879 19770 2175
rect 19200 1841 19262 1879
rect 19698 1841 19770 1879
rect 19950 2201 20250 2399
rect 19950 2149 20179 2201
rect 20231 2149 20250 2201
rect 19950 1941 20250 2149
rect 19950 1889 20179 1941
rect 20231 1889 20250 1941
rect 19950 1855 20250 1889
rect 20290 5986 20590 6150
rect 20290 5934 20309 5986
rect 20361 5934 20590 5986
rect 20290 5726 20590 5934
rect 20290 5674 20309 5726
rect 20361 5674 20590 5726
rect 20290 5476 20590 5674
rect 20290 5424 20309 5476
rect 20361 5424 20590 5476
rect 20290 5216 20590 5424
rect 20290 5164 20309 5216
rect 20361 5164 20590 5216
rect 20290 4956 20590 5164
rect 20290 4904 20309 4956
rect 20361 4904 20590 4956
rect 20290 4706 20590 4904
rect 20290 4654 20309 4706
rect 20361 4654 20590 4706
rect 20290 4446 20590 4654
rect 20290 4394 20309 4446
rect 20361 4394 20590 4446
rect 20290 4196 20590 4394
rect 20290 4144 20309 4196
rect 20361 4160 20590 4196
rect 20700 5476 21000 5490
rect 20700 5424 20929 5476
rect 20981 5424 21000 5476
rect 20700 5216 21000 5424
rect 20700 5164 20929 5216
rect 20981 5164 21000 5216
rect 20700 4966 21000 5164
rect 20700 4914 20929 4966
rect 20981 4914 21000 4966
rect 20700 4706 21000 4914
rect 20700 4654 20929 4706
rect 20981 4654 21000 4706
rect 20700 4446 21000 4654
rect 20700 4394 20929 4446
rect 20981 4394 21000 4446
rect 20700 4196 21000 4394
rect 21040 5346 21340 6300
rect 21040 5294 21059 5346
rect 21111 5294 21340 5346
rect 21040 5091 21340 5294
rect 21040 5039 21059 5091
rect 21111 5039 21340 5091
rect 21040 4836 21340 5039
rect 21040 4784 21059 4836
rect 21111 4784 21340 4836
rect 21040 4576 21340 4784
rect 21040 4524 21059 4576
rect 21111 4524 21340 4576
rect 21040 4316 21340 4524
rect 21040 4264 21059 4316
rect 21111 4264 21340 4316
rect 21040 4260 21340 4264
rect 21040 4250 21130 4260
rect 20700 4160 20929 4196
rect 20361 4144 20929 4160
rect 20981 4144 21000 4196
rect 20290 3871 21000 4144
rect 20290 3861 20929 3871
rect 20290 3809 20309 3861
rect 20361 3855 20929 3861
rect 20361 3809 20590 3855
rect 20290 3611 20590 3809
rect 20290 3559 20309 3611
rect 20361 3559 20590 3611
rect 20290 3351 20590 3559
rect 20290 3299 20309 3351
rect 20361 3299 20590 3351
rect 20290 3101 20590 3299
rect 20290 3049 20309 3101
rect 20361 3049 20590 3101
rect 20290 2841 20590 3049
rect 20290 2789 20309 2841
rect 20361 2789 20590 2841
rect 20290 2581 20590 2789
rect 20290 2529 20309 2581
rect 20361 2529 20590 2581
rect 20290 2331 20590 2529
rect 20700 3819 20929 3855
rect 20981 3819 21000 3871
rect 20700 3621 21000 3819
rect 20700 3569 20929 3621
rect 20981 3569 21000 3621
rect 20700 3361 21000 3569
rect 20700 3309 20929 3361
rect 20981 3309 21000 3361
rect 20700 3101 21000 3309
rect 20700 3049 20929 3101
rect 20981 3049 21000 3101
rect 20700 2851 21000 3049
rect 20700 2799 20929 2851
rect 20981 2799 21000 2851
rect 20700 2591 21000 2799
rect 20700 2539 20929 2591
rect 20981 2539 21000 2591
rect 20700 2520 21000 2539
rect 21040 3751 21340 3765
rect 21040 3699 21059 3751
rect 21111 3699 21340 3751
rect 21040 3491 21340 3699
rect 21040 3439 21059 3491
rect 21111 3439 21340 3491
rect 21040 3231 21340 3439
rect 21040 3179 21059 3231
rect 21111 3179 21340 3231
rect 21040 2976 21340 3179
rect 21040 2924 21059 2976
rect 21111 2924 21340 2976
rect 21040 2721 21340 2924
rect 21040 2669 21059 2721
rect 21111 2669 21340 2721
rect 20290 2279 20309 2331
rect 20361 2279 20590 2331
rect 20290 2071 20590 2279
rect 20290 2019 20309 2071
rect 20361 2019 20590 2071
rect 20290 1855 20590 2019
rect 19200 1805 19770 1841
rect 18500 1629 18514 1681
rect 18566 1629 19100 1681
rect 18500 1421 19100 1629
rect 18500 1369 18514 1421
rect 18566 1369 19100 1421
rect 18500 1171 19100 1369
rect 21040 1310 21340 2669
rect 18500 1119 18514 1171
rect 18566 1119 19100 1171
rect 18500 911 19100 1119
rect 18500 859 18514 911
rect 18566 859 19100 911
rect 19240 1249 21340 1310
rect 19240 941 19245 1249
rect 19745 941 21340 1249
rect 19240 880 21340 941
rect 18500 661 19100 859
rect 18500 609 18514 661
rect 18566 609 19100 661
rect 17190 349 17724 401
rect 17776 349 17790 401
rect 17190 285 17790 349
rect 18500 401 19100 609
rect 18500 349 18514 401
rect 18566 349 19100 401
rect 18500 285 19100 349
rect 16970 -132 18090 285
rect 16970 -184 17414 -132
rect 17466 -137 18009 -132
rect 17466 -184 17799 -137
rect 16970 -189 17799 -184
rect 17851 -184 18009 -137
rect 18061 -184 18090 -132
rect 17851 -189 18090 -184
rect 16970 -252 18090 -189
rect 16970 -304 17081 -252
rect 17133 -304 17271 -252
rect 17323 -304 17466 -252
rect 17518 -304 17656 -252
rect 17708 -304 17851 -252
rect 17903 -304 18090 -252
rect 16970 -315 18090 -304
rect 18195 -40 20515 285
rect 18195 -240 19315 -40
rect 18195 -252 19320 -240
rect 18195 -304 18386 -252
rect 18438 -304 18581 -252
rect 18633 -304 18771 -252
rect 18823 -304 18966 -252
rect 19018 -304 19156 -252
rect 19208 -304 19320 -252
rect 18195 -315 19320 -304
rect 16965 -377 19765 -365
rect 16965 -429 16981 -377
rect 17033 -429 17176 -377
rect 17228 -429 17371 -377
rect 17423 -429 17561 -377
rect 17613 -429 17751 -377
rect 17803 -429 17946 -377
rect 17998 -429 18291 -377
rect 18343 -429 18486 -377
rect 18538 -429 18676 -377
rect 18728 -429 18866 -377
rect 18918 -429 19061 -377
rect 19113 -397 19256 -377
rect 19308 -397 19765 -377
rect 19113 -429 19252 -397
rect 16965 -933 19252 -429
rect 19708 -933 19765 -397
rect 16965 -965 19765 -933
<< via2 >>
rect 17469 7179 17525 7235
rect 17549 7179 17605 7235
rect 17629 7179 17685 7235
rect 18124 7179 18180 7235
rect 18204 7179 18260 7235
rect 18284 7179 18340 7235
rect 18769 7179 18825 7235
rect 18849 7179 18905 7235
rect 18929 7179 18985 7235
rect 19992 6064 20179 6098
rect 20179 6064 20208 6098
rect 19992 5962 20208 6064
rect 19252 1879 19262 2175
rect 19262 1879 19698 2175
rect 19698 1879 19708 2175
rect 19252 -429 19256 -397
rect 19256 -429 19308 -397
rect 19308 -429 19708 -397
rect 19252 -933 19708 -429
<< metal3 >>
rect 17440 7235 20250 7275
rect 17440 7179 17469 7235
rect 17525 7179 17549 7235
rect 17605 7179 17629 7235
rect 17685 7179 18124 7235
rect 18180 7179 18204 7235
rect 18260 7179 18284 7235
rect 18340 7179 18769 7235
rect 18825 7179 18849 7235
rect 18905 7179 18929 7235
rect 18985 7179 20250 7235
rect 17440 7140 20250 7179
rect 19950 6098 20250 7140
rect 19950 5962 19992 6098
rect 20208 5962 20250 6098
rect 19950 5905 20250 5962
rect 19200 2175 19770 2255
rect 19200 1879 19252 2175
rect 19708 1879 19770 2175
rect 19200 1805 19770 1879
rect 19200 -397 19765 1805
rect 19200 -933 19252 -397
rect 19708 -933 19765 -397
rect 19200 -965 19765 -933
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM1
timestamp 1663011646
transform 0 1 20269 -1 0 2877
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM2
timestamp 1663011646
transform 0 1 18069 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM3
timestamp 1663011646
transform 0 1 18719 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM29
timestamp 1663011646
transform 0 1 20269 -1 0 5127
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4  XM30
timestamp 1663011646
transform 0 1 21019 -1 0 3207
box -807 -319 807 319
use sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4  XM31
timestamp 1663011646
transform 0 1 21019 -1 0 4807
box -807 -319 807 319
use sky130_fd_pr__pfet_01v8_lvt_D3M934  XM36
timestamp 1663011646
transform 0 1 17419 -1 0 6117
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_lvt_D3Z634  XM37
timestamp 1663011646
transform 0 1 17819 -1 0 2297
box -2087 -319 2087 319
use sky130_fd_pr__pfet_01v8_lvt_D3Z634  XM38
timestamp 1663011646
transform 0 1 18469 -1 0 2297
box -2087 -319 2087 319
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM39
timestamp 1663011646
transform 1 0 17493 0 1 -340
box -637 -300 637 300
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM40
timestamp 1663011646
transform -1 0 18797 0 -1 -340
box -637 -300 637 300
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR19
timestamp 1663011646
transform 1 0 19491 0 1 5548
box -441 -1348 441 1348
use sky130_fd_pr__res_high_po_2p85_MM89SS  XR20
timestamp 1663011646
transform 1 0 19491 0 1 2448
box -441 -1728 441 1728
<< labels >>
rlabel metal1 s 20820 5520 21340 5580 4 AMP
port 1 nsew
rlabel metal1 s 21020 2435 21340 2495 4 VOP
port 2 nsew
rlabel metal3 s 18360 7140 18750 7275 4 VDD
port 3 nsew
rlabel metal2 s 19060 -40 20515 285 4 BIASOUT
port 4 nsew
rlabel locali s 18970 6975 20025 7020 4 PSUB
port 5 nsew
rlabel metal1 s 17220 7150 20470 7220 4 BIAS2V
port 6 nsew
rlabel metal1 s 17100 4310 18020 4370 4 VCTRL
port 7 nsew
rlabel metal2 s 16965 -965 19230 -430 4 GND
port 8 nsew
rlabel locali s 19070 -100 19115 790 4 SUB
port 9 nsew
<< end >>
