magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -812 -284 812 284
<< pmoslvt >>
rect -616 -136 -416 64
rect -358 -136 -158 64
rect -100 -136 100 64
rect 158 -136 358 64
rect 416 -136 616 64
<< pdiff >>
rect -674 49 -616 64
rect -674 15 -662 49
rect -628 15 -616 49
rect -674 -19 -616 15
rect -674 -53 -662 -19
rect -628 -53 -616 -19
rect -674 -87 -616 -53
rect -674 -121 -662 -87
rect -628 -121 -616 -87
rect -674 -136 -616 -121
rect -416 49 -358 64
rect -416 15 -404 49
rect -370 15 -358 49
rect -416 -19 -358 15
rect -416 -53 -404 -19
rect -370 -53 -358 -19
rect -416 -87 -358 -53
rect -416 -121 -404 -87
rect -370 -121 -358 -87
rect -416 -136 -358 -121
rect -158 49 -100 64
rect -158 15 -146 49
rect -112 15 -100 49
rect -158 -19 -100 15
rect -158 -53 -146 -19
rect -112 -53 -100 -19
rect -158 -87 -100 -53
rect -158 -121 -146 -87
rect -112 -121 -100 -87
rect -158 -136 -100 -121
rect 100 49 158 64
rect 100 15 112 49
rect 146 15 158 49
rect 100 -19 158 15
rect 100 -53 112 -19
rect 146 -53 158 -19
rect 100 -87 158 -53
rect 100 -121 112 -87
rect 146 -121 158 -87
rect 100 -136 158 -121
rect 358 49 416 64
rect 358 15 370 49
rect 404 15 416 49
rect 358 -19 416 15
rect 358 -53 370 -19
rect 404 -53 416 -19
rect 358 -87 416 -53
rect 358 -121 370 -87
rect 404 -121 416 -87
rect 358 -136 416 -121
rect 616 49 674 64
rect 616 15 628 49
rect 662 15 674 49
rect 616 -19 674 15
rect 616 -53 628 -19
rect 662 -53 674 -19
rect 616 -87 674 -53
rect 616 -121 628 -87
rect 662 -121 674 -87
rect 616 -136 674 -121
<< pdiffc >>
rect -662 15 -628 49
rect -662 -53 -628 -19
rect -662 -121 -628 -87
rect -404 15 -370 49
rect -404 -53 -370 -19
rect -404 -121 -370 -87
rect -146 15 -112 49
rect -146 -53 -112 -19
rect -146 -121 -112 -87
rect 112 15 146 49
rect 112 -53 146 -19
rect 112 -121 146 -87
rect 370 15 404 49
rect 370 -53 404 -19
rect 370 -121 404 -87
rect 628 15 662 49
rect 628 -53 662 -19
rect 628 -121 662 -87
<< nsubdiff >>
rect -776 214 776 248
rect -776 119 -742 214
rect -776 51 -742 85
rect 742 119 776 214
rect -776 -17 -742 17
rect -776 -85 -742 -51
rect -776 -214 -742 -119
rect 742 51 776 85
rect 742 -17 776 17
rect 742 -85 776 -51
rect 742 -214 776 -119
rect -776 -248 776 -214
<< nsubdiffcont >>
rect -776 85 -742 119
rect 742 85 776 119
rect -776 17 -742 51
rect -776 -51 -742 -17
rect -776 -119 -742 -85
rect 742 17 776 51
rect 742 -51 776 -17
rect 742 -119 776 -85
<< poly >>
rect -616 145 -416 161
rect -616 111 -567 145
rect -533 111 -499 145
rect -465 111 -416 145
rect -616 64 -416 111
rect -358 145 -158 161
rect -358 111 -309 145
rect -275 111 -241 145
rect -207 111 -158 145
rect -358 64 -158 111
rect -100 145 100 161
rect -100 111 -51 145
rect -17 111 17 145
rect 51 111 100 145
rect -100 64 100 111
rect 158 145 358 161
rect 158 111 207 145
rect 241 111 275 145
rect 309 111 358 145
rect 158 64 358 111
rect 416 145 616 161
rect 416 111 465 145
rect 499 111 533 145
rect 567 111 616 145
rect 416 64 616 111
rect -616 -162 -416 -136
rect -358 -162 -158 -136
rect -100 -162 100 -136
rect 158 -162 358 -136
rect 416 -162 616 -136
<< polycont >>
rect -567 111 -533 145
rect -499 111 -465 145
rect -309 111 -275 145
rect -241 111 -207 145
rect -51 111 -17 145
rect 17 111 51 145
rect 207 111 241 145
rect 275 111 309 145
rect 465 111 499 145
rect 533 111 567 145
<< locali >>
rect -776 214 776 248
rect -776 119 -742 214
rect -616 111 -569 145
rect -533 111 -499 145
rect -463 111 -416 145
rect -358 111 -311 145
rect -275 111 -241 145
rect -205 111 -158 145
rect -100 111 -53 145
rect -17 111 17 145
rect 53 111 100 145
rect 158 111 205 145
rect 241 111 275 145
rect 311 111 358 145
rect 416 111 463 145
rect 499 111 533 145
rect 569 111 616 145
rect 742 119 776 214
rect -776 51 -742 85
rect -776 -17 -742 17
rect -776 -85 -742 -51
rect -776 -214 -742 -119
rect -662 49 -628 68
rect -662 -19 -628 -17
rect -662 -55 -628 -53
rect -662 -140 -628 -121
rect -404 49 -370 68
rect -404 -19 -370 -17
rect -404 -55 -370 -53
rect -404 -140 -370 -121
rect -146 49 -112 68
rect -146 -19 -112 -17
rect -146 -55 -112 -53
rect -146 -140 -112 -121
rect 112 49 146 68
rect 112 -19 146 -17
rect 112 -55 146 -53
rect 112 -140 146 -121
rect 370 49 404 68
rect 370 -19 404 -17
rect 370 -55 404 -53
rect 370 -140 404 -121
rect 628 49 662 68
rect 628 -19 662 -17
rect 628 -55 662 -53
rect 628 -140 662 -121
rect 742 51 776 85
rect 742 -17 776 17
rect 742 -85 776 -51
rect 742 -214 776 -119
rect -776 -248 776 -214
<< viali >>
rect -569 111 -567 145
rect -567 111 -535 145
rect -497 111 -465 145
rect -465 111 -463 145
rect -311 111 -309 145
rect -309 111 -277 145
rect -239 111 -207 145
rect -207 111 -205 145
rect -53 111 -51 145
rect -51 111 -19 145
rect 19 111 51 145
rect 51 111 53 145
rect 205 111 207 145
rect 207 111 239 145
rect 277 111 309 145
rect 309 111 311 145
rect 463 111 465 145
rect 465 111 497 145
rect 535 111 567 145
rect 567 111 569 145
rect -662 15 -628 17
rect -662 -17 -628 15
rect -662 -87 -628 -55
rect -662 -89 -628 -87
rect -404 15 -370 17
rect -404 -17 -370 15
rect -404 -87 -370 -55
rect -404 -89 -370 -87
rect -146 15 -112 17
rect -146 -17 -112 15
rect -146 -87 -112 -55
rect -146 -89 -112 -87
rect 112 15 146 17
rect 112 -17 146 15
rect 112 -87 146 -55
rect 112 -89 146 -87
rect 370 15 404 17
rect 370 -17 404 15
rect 370 -87 404 -55
rect 370 -89 404 -87
rect 628 15 662 17
rect 628 -17 662 15
rect 628 -87 662 -55
rect 628 -89 662 -87
<< metal1 >>
rect -612 145 -420 151
rect -612 111 -569 145
rect -535 111 -497 145
rect -463 111 -420 145
rect -612 105 -420 111
rect -354 145 -162 151
rect -354 111 -311 145
rect -277 111 -239 145
rect -205 111 -162 145
rect -354 105 -162 111
rect -96 145 96 151
rect -96 111 -53 145
rect -19 111 19 145
rect 53 111 96 145
rect -96 105 96 111
rect 162 145 354 151
rect 162 111 205 145
rect 239 111 277 145
rect 311 111 354 145
rect 162 105 354 111
rect 420 145 612 151
rect 420 111 463 145
rect 497 111 535 145
rect 569 111 612 145
rect 420 105 612 111
rect -668 17 -622 64
rect -668 -17 -662 17
rect -628 -17 -622 17
rect -668 -55 -622 -17
rect -668 -89 -662 -55
rect -628 -89 -622 -55
rect -668 -136 -622 -89
rect -410 17 -364 64
rect -410 -17 -404 17
rect -370 -17 -364 17
rect -410 -55 -364 -17
rect -410 -89 -404 -55
rect -370 -89 -364 -55
rect -410 -136 -364 -89
rect -152 17 -106 64
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -55 -106 -17
rect -152 -89 -146 -55
rect -112 -89 -106 -55
rect -152 -136 -106 -89
rect 106 17 152 64
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -55 152 -17
rect 106 -89 112 -55
rect 146 -89 152 -55
rect 106 -136 152 -89
rect 364 17 410 64
rect 364 -17 370 17
rect 404 -17 410 17
rect 364 -55 410 -17
rect 364 -89 370 -55
rect 404 -89 410 -55
rect 364 -136 410 -89
rect 622 17 668 64
rect 622 -17 628 17
rect 662 -17 668 17
rect 622 -55 668 -17
rect 622 -89 628 -55
rect 662 -89 668 -55
rect 622 -136 668 -89
<< properties >>
string FIXED_BBOX -759 -231 759 231
<< end >>
