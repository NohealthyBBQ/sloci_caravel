magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 5840 10060 6580 10100
rect 7190 10060 7410 10100
rect 7990 10060 8210 10100
rect 8790 10060 9010 10100
rect 5840 9550 6590 9590
rect 7190 9540 7410 9580
rect 7990 9540 8210 9580
rect 8790 9540 9010 9580
<< metal1 >>
rect 5160 9974 5740 10040
rect 5160 9666 5200 9974
rect 5700 9666 5740 9974
rect 5160 9600 5740 9666
rect 6570 10010 6640 10130
rect 7370 10010 7440 10130
rect 8170 10010 8240 10130
rect 8970 10010 9040 10130
rect 6570 9950 6980 10010
rect 7370 9950 7780 10010
rect 8170 9950 8580 10010
rect 8970 9950 9380 10010
rect 6570 9690 6640 9950
rect 6670 9906 6750 9920
rect 6670 9854 6684 9906
rect 6736 9854 6750 9906
rect 6670 9840 6750 9854
rect 6680 9720 6730 9840
rect 6780 9800 6830 9920
rect 6860 9906 6940 9920
rect 6860 9854 6874 9906
rect 6926 9854 6940 9906
rect 6860 9840 6940 9854
rect 6760 9786 6840 9800
rect 6760 9734 6774 9786
rect 6826 9734 6840 9786
rect 6760 9720 6840 9734
rect 6870 9720 6930 9840
rect 6970 9810 7030 9920
rect 7060 9906 7140 9920
rect 7060 9854 7074 9906
rect 7126 9854 7140 9906
rect 7060 9840 7140 9854
rect 7060 9830 7120 9840
rect 6960 9800 7030 9810
rect 6960 9786 7040 9800
rect 6960 9734 6974 9786
rect 7026 9734 7040 9786
rect 6960 9720 7040 9734
rect 7070 9720 7120 9830
rect 7370 9690 7440 9950
rect 7470 9906 7550 9920
rect 7470 9854 7484 9906
rect 7536 9854 7550 9906
rect 7470 9840 7550 9854
rect 7480 9720 7530 9840
rect 7580 9800 7630 9920
rect 7660 9906 7740 9920
rect 7660 9854 7674 9906
rect 7726 9854 7740 9906
rect 7660 9840 7740 9854
rect 7560 9786 7640 9800
rect 7560 9734 7574 9786
rect 7626 9734 7640 9786
rect 7560 9720 7640 9734
rect 7670 9720 7730 9840
rect 7770 9810 7830 9920
rect 7860 9906 7940 9920
rect 7860 9854 7874 9906
rect 7926 9854 7940 9906
rect 7860 9840 7940 9854
rect 7860 9830 7920 9840
rect 7760 9800 7830 9810
rect 7760 9786 7840 9800
rect 7760 9734 7774 9786
rect 7826 9734 7840 9786
rect 7760 9720 7840 9734
rect 7868 9720 7920 9830
rect 8170 9690 8240 9950
rect 8270 9906 8350 9920
rect 8270 9854 8284 9906
rect 8336 9854 8350 9906
rect 8270 9840 8350 9854
rect 8280 9720 8330 9840
rect 8380 9800 8430 9920
rect 8460 9906 8540 9920
rect 8460 9854 8474 9906
rect 8526 9854 8540 9906
rect 8460 9840 8540 9854
rect 8360 9786 8440 9800
rect 8360 9734 8374 9786
rect 8426 9734 8440 9786
rect 8360 9720 8440 9734
rect 8470 9720 8530 9840
rect 8570 9810 8630 9920
rect 8660 9906 8740 9920
rect 8660 9854 8674 9906
rect 8726 9854 8740 9906
rect 8660 9840 8740 9854
rect 8660 9830 8720 9840
rect 8560 9800 8630 9810
rect 8560 9786 8640 9800
rect 8560 9734 8574 9786
rect 8626 9734 8640 9786
rect 8560 9720 8640 9734
rect 8668 9720 8720 9830
rect 8970 9690 9040 9950
rect 9070 9906 9150 9920
rect 9070 9854 9084 9906
rect 9136 9854 9150 9906
rect 9070 9840 9150 9854
rect 9080 9720 9130 9840
rect 9180 9800 9230 9920
rect 9260 9906 9340 9920
rect 9260 9854 9274 9906
rect 9326 9854 9340 9906
rect 9260 9840 9340 9854
rect 9160 9786 9240 9800
rect 9160 9734 9174 9786
rect 9226 9734 9240 9786
rect 9160 9720 9240 9734
rect 9270 9720 9330 9840
rect 9370 9810 9430 9920
rect 9460 9906 9540 9920
rect 9460 9854 9474 9906
rect 9526 9854 9540 9906
rect 9460 9840 9540 9854
rect 9460 9830 9520 9840
rect 9360 9800 9430 9810
rect 9360 9786 9440 9800
rect 9360 9734 9374 9786
rect 9426 9734 9440 9786
rect 9360 9720 9440 9734
rect 9468 9720 9520 9830
rect 6570 9640 7080 9690
rect 7370 9640 7880 9690
rect 8170 9640 8680 9690
rect 8970 9640 9480 9690
rect 5100 1188 5780 1240
rect 5100 752 5158 1188
rect 5722 752 5780 1188
rect 5100 700 5780 752
<< via1 >>
rect 5200 9666 5700 9974
rect 6684 9854 6736 9906
rect 6874 9854 6926 9906
rect 6774 9734 6826 9786
rect 7074 9854 7126 9906
rect 6974 9734 7026 9786
rect 7484 9854 7536 9906
rect 7674 9854 7726 9906
rect 7574 9734 7626 9786
rect 7874 9854 7926 9906
rect 7774 9734 7826 9786
rect 8284 9854 8336 9906
rect 8474 9854 8526 9906
rect 8374 9734 8426 9786
rect 8674 9854 8726 9906
rect 8574 9734 8626 9786
rect 9084 9854 9136 9906
rect 9274 9854 9326 9906
rect 9174 9734 9226 9786
rect 9474 9854 9526 9906
rect 9374 9734 9426 9786
rect 5158 752 5722 1188
<< metal2 >>
rect 7670 10040 7870 10060
rect 8470 10040 8670 10060
rect 9270 10040 9470 10060
rect 5160 9988 9540 10040
rect 5160 9974 6092 9988
rect 5160 9666 5200 9974
rect 5700 9692 6092 9974
rect 6388 9906 9540 9988
rect 6388 9854 6684 9906
rect 6736 9854 6874 9906
rect 6926 9854 7074 9906
rect 7126 9854 7484 9906
rect 7536 9854 7674 9906
rect 7726 9854 7874 9906
rect 7926 9854 8284 9906
rect 8336 9854 8474 9906
rect 8526 9854 8674 9906
rect 8726 9854 9084 9906
rect 9136 9854 9274 9906
rect 9326 9854 9474 9906
rect 9526 9854 9540 9906
rect 6388 9840 9540 9854
rect 6388 9692 6440 9840
rect 5700 9666 6440 9692
rect 5160 9640 6440 9666
rect 6540 9786 9570 9800
rect 6540 9734 6774 9786
rect 6826 9734 6974 9786
rect 7026 9734 7574 9786
rect 7626 9734 7774 9786
rect 7826 9734 8374 9786
rect 8426 9734 8574 9786
rect 8626 9734 9174 9786
rect 9226 9734 9374 9786
rect 9426 9734 9570 9786
rect 5160 9600 5740 9640
rect 6540 9510 9570 9734
rect 6540 9360 6830 9510
rect 5000 9070 6830 9360
rect 5000 1198 5780 1240
rect 5000 1188 5172 1198
rect 5708 1188 5780 1198
rect 5000 752 5158 1188
rect 5722 752 5780 1188
rect 5000 742 5172 752
rect 5708 742 5780 752
rect 5000 600 5780 742
<< via2 >>
rect 6092 9692 6388 9988
rect 5172 1188 5708 1198
rect 5172 752 5708 1188
rect 5172 742 5708 752
<< metal3 >>
rect 6040 9992 6440 10040
rect 6040 9688 6088 9992
rect 6392 9688 6440 9992
rect 6040 9640 6440 9688
rect 5100 1198 6040 1240
rect 5100 742 5172 1198
rect 5708 742 6040 1198
rect 5100 700 6040 742
<< via3 >>
rect 6088 9988 6392 9992
rect 6088 9692 6092 9988
rect 6092 9692 6388 9988
rect 6388 9692 6392 9988
rect 6088 9688 6392 9692
<< metal4 >>
rect 6040 9992 6440 10040
rect 6040 9688 6088 9992
rect 6392 9688 6440 9992
rect 6040 6420 6440 9688
rect 6040 590 6430 1670
use sky130_fd_pr__cap_mim_m3_1_4RCNTW  XC1
timestamp 1663011646
transform 1 0 8050 0 1 3700
box -2150 -3100 2149 3100
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM25
timestamp 1663011646
transform 1 0 8499 0 -1 9820
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM26
timestamp 1663011646
transform 1 0 9299 0 -1 9820
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM27
timestamp 1663011646
transform 1 0 7699 0 -1 9820
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM28
timestamp 1663011646
transform 1 0 6899 0 -1 9820
box -349 -300 349 300
use sky130_fd_pr__res_high_po_2p85_MXEQGY  XR18
timestamp 1663011646
transform 1 0 5451 0 1 5398
box -441 -4788 441 4788
<< labels >>
rlabel metal2 s 5000 600 5140 1240 4 GND
port 1 nsew
rlabel metal1 s 6570 9950 6640 10130 4 IN1
port 2 nsew
rlabel metal2 s 5000 9070 6830 9360 4 VDD
port 3 nsew
rlabel metal1 s 7370 9640 7440 10130 4 IN2
port 4 nsew
rlabel metal1 s 8170 9640 8240 10130 4 IN3
port 5 nsew
rlabel metal1 s 8970 9640 9040 10130 4 IN4
port 6 nsew
rlabel metal4 s 6040 590 6430 1670 4 AMP
port 7 nsew
rlabel locali s 5840 10060 6580 10100 4 SUB
port 8 nsew
<< end >>
