magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -971 -857 971 795
<< nmoslvt >>
rect -887 -831 -487 769
rect -429 -831 -29 769
rect 29 -831 429 769
rect 487 -831 887 769
<< ndiff >>
rect -945 734 -887 769
rect -945 700 -933 734
rect -899 700 -887 734
rect -945 666 -887 700
rect -945 632 -933 666
rect -899 632 -887 666
rect -945 598 -887 632
rect -945 564 -933 598
rect -899 564 -887 598
rect -945 530 -887 564
rect -945 496 -933 530
rect -899 496 -887 530
rect -945 462 -887 496
rect -945 428 -933 462
rect -899 428 -887 462
rect -945 394 -887 428
rect -945 360 -933 394
rect -899 360 -887 394
rect -945 326 -887 360
rect -945 292 -933 326
rect -899 292 -887 326
rect -945 258 -887 292
rect -945 224 -933 258
rect -899 224 -887 258
rect -945 190 -887 224
rect -945 156 -933 190
rect -899 156 -887 190
rect -945 122 -887 156
rect -945 88 -933 122
rect -899 88 -887 122
rect -945 54 -887 88
rect -945 20 -933 54
rect -899 20 -887 54
rect -945 -14 -887 20
rect -945 -48 -933 -14
rect -899 -48 -887 -14
rect -945 -82 -887 -48
rect -945 -116 -933 -82
rect -899 -116 -887 -82
rect -945 -150 -887 -116
rect -945 -184 -933 -150
rect -899 -184 -887 -150
rect -945 -218 -887 -184
rect -945 -252 -933 -218
rect -899 -252 -887 -218
rect -945 -286 -887 -252
rect -945 -320 -933 -286
rect -899 -320 -887 -286
rect -945 -354 -887 -320
rect -945 -388 -933 -354
rect -899 -388 -887 -354
rect -945 -422 -887 -388
rect -945 -456 -933 -422
rect -899 -456 -887 -422
rect -945 -490 -887 -456
rect -945 -524 -933 -490
rect -899 -524 -887 -490
rect -945 -558 -887 -524
rect -945 -592 -933 -558
rect -899 -592 -887 -558
rect -945 -626 -887 -592
rect -945 -660 -933 -626
rect -899 -660 -887 -626
rect -945 -694 -887 -660
rect -945 -728 -933 -694
rect -899 -728 -887 -694
rect -945 -762 -887 -728
rect -945 -796 -933 -762
rect -899 -796 -887 -762
rect -945 -831 -887 -796
rect -487 734 -429 769
rect -487 700 -475 734
rect -441 700 -429 734
rect -487 666 -429 700
rect -487 632 -475 666
rect -441 632 -429 666
rect -487 598 -429 632
rect -487 564 -475 598
rect -441 564 -429 598
rect -487 530 -429 564
rect -487 496 -475 530
rect -441 496 -429 530
rect -487 462 -429 496
rect -487 428 -475 462
rect -441 428 -429 462
rect -487 394 -429 428
rect -487 360 -475 394
rect -441 360 -429 394
rect -487 326 -429 360
rect -487 292 -475 326
rect -441 292 -429 326
rect -487 258 -429 292
rect -487 224 -475 258
rect -441 224 -429 258
rect -487 190 -429 224
rect -487 156 -475 190
rect -441 156 -429 190
rect -487 122 -429 156
rect -487 88 -475 122
rect -441 88 -429 122
rect -487 54 -429 88
rect -487 20 -475 54
rect -441 20 -429 54
rect -487 -14 -429 20
rect -487 -48 -475 -14
rect -441 -48 -429 -14
rect -487 -82 -429 -48
rect -487 -116 -475 -82
rect -441 -116 -429 -82
rect -487 -150 -429 -116
rect -487 -184 -475 -150
rect -441 -184 -429 -150
rect -487 -218 -429 -184
rect -487 -252 -475 -218
rect -441 -252 -429 -218
rect -487 -286 -429 -252
rect -487 -320 -475 -286
rect -441 -320 -429 -286
rect -487 -354 -429 -320
rect -487 -388 -475 -354
rect -441 -388 -429 -354
rect -487 -422 -429 -388
rect -487 -456 -475 -422
rect -441 -456 -429 -422
rect -487 -490 -429 -456
rect -487 -524 -475 -490
rect -441 -524 -429 -490
rect -487 -558 -429 -524
rect -487 -592 -475 -558
rect -441 -592 -429 -558
rect -487 -626 -429 -592
rect -487 -660 -475 -626
rect -441 -660 -429 -626
rect -487 -694 -429 -660
rect -487 -728 -475 -694
rect -441 -728 -429 -694
rect -487 -762 -429 -728
rect -487 -796 -475 -762
rect -441 -796 -429 -762
rect -487 -831 -429 -796
rect -29 734 29 769
rect -29 700 -17 734
rect 17 700 29 734
rect -29 666 29 700
rect -29 632 -17 666
rect 17 632 29 666
rect -29 598 29 632
rect -29 564 -17 598
rect 17 564 29 598
rect -29 530 29 564
rect -29 496 -17 530
rect 17 496 29 530
rect -29 462 29 496
rect -29 428 -17 462
rect 17 428 29 462
rect -29 394 29 428
rect -29 360 -17 394
rect 17 360 29 394
rect -29 326 29 360
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -422 29 -388
rect -29 -456 -17 -422
rect 17 -456 29 -422
rect -29 -490 29 -456
rect -29 -524 -17 -490
rect 17 -524 29 -490
rect -29 -558 29 -524
rect -29 -592 -17 -558
rect 17 -592 29 -558
rect -29 -626 29 -592
rect -29 -660 -17 -626
rect 17 -660 29 -626
rect -29 -694 29 -660
rect -29 -728 -17 -694
rect 17 -728 29 -694
rect -29 -762 29 -728
rect -29 -796 -17 -762
rect 17 -796 29 -762
rect -29 -831 29 -796
rect 429 734 487 769
rect 429 700 441 734
rect 475 700 487 734
rect 429 666 487 700
rect 429 632 441 666
rect 475 632 487 666
rect 429 598 487 632
rect 429 564 441 598
rect 475 564 487 598
rect 429 530 487 564
rect 429 496 441 530
rect 475 496 487 530
rect 429 462 487 496
rect 429 428 441 462
rect 475 428 487 462
rect 429 394 487 428
rect 429 360 441 394
rect 475 360 487 394
rect 429 326 487 360
rect 429 292 441 326
rect 475 292 487 326
rect 429 258 487 292
rect 429 224 441 258
rect 475 224 487 258
rect 429 190 487 224
rect 429 156 441 190
rect 475 156 487 190
rect 429 122 487 156
rect 429 88 441 122
rect 475 88 487 122
rect 429 54 487 88
rect 429 20 441 54
rect 475 20 487 54
rect 429 -14 487 20
rect 429 -48 441 -14
rect 475 -48 487 -14
rect 429 -82 487 -48
rect 429 -116 441 -82
rect 475 -116 487 -82
rect 429 -150 487 -116
rect 429 -184 441 -150
rect 475 -184 487 -150
rect 429 -218 487 -184
rect 429 -252 441 -218
rect 475 -252 487 -218
rect 429 -286 487 -252
rect 429 -320 441 -286
rect 475 -320 487 -286
rect 429 -354 487 -320
rect 429 -388 441 -354
rect 475 -388 487 -354
rect 429 -422 487 -388
rect 429 -456 441 -422
rect 475 -456 487 -422
rect 429 -490 487 -456
rect 429 -524 441 -490
rect 475 -524 487 -490
rect 429 -558 487 -524
rect 429 -592 441 -558
rect 475 -592 487 -558
rect 429 -626 487 -592
rect 429 -660 441 -626
rect 475 -660 487 -626
rect 429 -694 487 -660
rect 429 -728 441 -694
rect 475 -728 487 -694
rect 429 -762 487 -728
rect 429 -796 441 -762
rect 475 -796 487 -762
rect 429 -831 487 -796
rect 887 734 945 769
rect 887 700 899 734
rect 933 700 945 734
rect 887 666 945 700
rect 887 632 899 666
rect 933 632 945 666
rect 887 598 945 632
rect 887 564 899 598
rect 933 564 945 598
rect 887 530 945 564
rect 887 496 899 530
rect 933 496 945 530
rect 887 462 945 496
rect 887 428 899 462
rect 933 428 945 462
rect 887 394 945 428
rect 887 360 899 394
rect 933 360 945 394
rect 887 326 945 360
rect 887 292 899 326
rect 933 292 945 326
rect 887 258 945 292
rect 887 224 899 258
rect 933 224 945 258
rect 887 190 945 224
rect 887 156 899 190
rect 933 156 945 190
rect 887 122 945 156
rect 887 88 899 122
rect 933 88 945 122
rect 887 54 945 88
rect 887 20 899 54
rect 933 20 945 54
rect 887 -14 945 20
rect 887 -48 899 -14
rect 933 -48 945 -14
rect 887 -82 945 -48
rect 887 -116 899 -82
rect 933 -116 945 -82
rect 887 -150 945 -116
rect 887 -184 899 -150
rect 933 -184 945 -150
rect 887 -218 945 -184
rect 887 -252 899 -218
rect 933 -252 945 -218
rect 887 -286 945 -252
rect 887 -320 899 -286
rect 933 -320 945 -286
rect 887 -354 945 -320
rect 887 -388 899 -354
rect 933 -388 945 -354
rect 887 -422 945 -388
rect 887 -456 899 -422
rect 933 -456 945 -422
rect 887 -490 945 -456
rect 887 -524 899 -490
rect 933 -524 945 -490
rect 887 -558 945 -524
rect 887 -592 899 -558
rect 933 -592 945 -558
rect 887 -626 945 -592
rect 887 -660 899 -626
rect 933 -660 945 -626
rect 887 -694 945 -660
rect 887 -728 899 -694
rect 933 -728 945 -694
rect 887 -762 945 -728
rect 887 -796 899 -762
rect 933 -796 945 -762
rect 887 -831 945 -796
<< ndiffc >>
rect -933 700 -899 734
rect -933 632 -899 666
rect -933 564 -899 598
rect -933 496 -899 530
rect -933 428 -899 462
rect -933 360 -899 394
rect -933 292 -899 326
rect -933 224 -899 258
rect -933 156 -899 190
rect -933 88 -899 122
rect -933 20 -899 54
rect -933 -48 -899 -14
rect -933 -116 -899 -82
rect -933 -184 -899 -150
rect -933 -252 -899 -218
rect -933 -320 -899 -286
rect -933 -388 -899 -354
rect -933 -456 -899 -422
rect -933 -524 -899 -490
rect -933 -592 -899 -558
rect -933 -660 -899 -626
rect -933 -728 -899 -694
rect -933 -796 -899 -762
rect -475 700 -441 734
rect -475 632 -441 666
rect -475 564 -441 598
rect -475 496 -441 530
rect -475 428 -441 462
rect -475 360 -441 394
rect -475 292 -441 326
rect -475 224 -441 258
rect -475 156 -441 190
rect -475 88 -441 122
rect -475 20 -441 54
rect -475 -48 -441 -14
rect -475 -116 -441 -82
rect -475 -184 -441 -150
rect -475 -252 -441 -218
rect -475 -320 -441 -286
rect -475 -388 -441 -354
rect -475 -456 -441 -422
rect -475 -524 -441 -490
rect -475 -592 -441 -558
rect -475 -660 -441 -626
rect -475 -728 -441 -694
rect -475 -796 -441 -762
rect -17 700 17 734
rect -17 632 17 666
rect -17 564 17 598
rect -17 496 17 530
rect -17 428 17 462
rect -17 360 17 394
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect -17 -456 17 -422
rect -17 -524 17 -490
rect -17 -592 17 -558
rect -17 -660 17 -626
rect -17 -728 17 -694
rect -17 -796 17 -762
rect 441 700 475 734
rect 441 632 475 666
rect 441 564 475 598
rect 441 496 475 530
rect 441 428 475 462
rect 441 360 475 394
rect 441 292 475 326
rect 441 224 475 258
rect 441 156 475 190
rect 441 88 475 122
rect 441 20 475 54
rect 441 -48 475 -14
rect 441 -116 475 -82
rect 441 -184 475 -150
rect 441 -252 475 -218
rect 441 -320 475 -286
rect 441 -388 475 -354
rect 441 -456 475 -422
rect 441 -524 475 -490
rect 441 -592 475 -558
rect 441 -660 475 -626
rect 441 -728 475 -694
rect 441 -796 475 -762
rect 899 700 933 734
rect 899 632 933 666
rect 899 564 933 598
rect 899 496 933 530
rect 899 428 933 462
rect 899 360 933 394
rect 899 292 933 326
rect 899 224 933 258
rect 899 156 933 190
rect 899 88 933 122
rect 899 20 933 54
rect 899 -48 933 -14
rect 899 -116 933 -82
rect 899 -184 933 -150
rect 899 -252 933 -218
rect 899 -320 933 -286
rect 899 -388 933 -354
rect 899 -456 933 -422
rect 899 -524 933 -490
rect 899 -592 933 -558
rect 899 -660 933 -626
rect 899 -728 933 -694
rect 899 -796 933 -762
<< poly >>
rect -887 841 -487 857
rect -887 807 -840 841
rect -806 807 -772 841
rect -738 807 -704 841
rect -670 807 -636 841
rect -602 807 -568 841
rect -534 807 -487 841
rect -887 769 -487 807
rect -429 841 -29 857
rect -429 807 -382 841
rect -348 807 -314 841
rect -280 807 -246 841
rect -212 807 -178 841
rect -144 807 -110 841
rect -76 807 -29 841
rect -429 769 -29 807
rect 29 841 429 857
rect 29 807 76 841
rect 110 807 144 841
rect 178 807 212 841
rect 246 807 280 841
rect 314 807 348 841
rect 382 807 429 841
rect 29 769 429 807
rect 487 841 887 857
rect 487 807 534 841
rect 568 807 602 841
rect 636 807 670 841
rect 704 807 738 841
rect 772 807 806 841
rect 840 807 887 841
rect 487 769 887 807
rect -887 -857 -487 -831
rect -429 -857 -29 -831
rect 29 -857 429 -831
rect 487 -857 887 -831
<< polycont >>
rect -840 807 -806 841
rect -772 807 -738 841
rect -704 807 -670 841
rect -636 807 -602 841
rect -568 807 -534 841
rect -382 807 -348 841
rect -314 807 -280 841
rect -246 807 -212 841
rect -178 807 -144 841
rect -110 807 -76 841
rect 76 807 110 841
rect 144 807 178 841
rect 212 807 246 841
rect 280 807 314 841
rect 348 807 382 841
rect 534 807 568 841
rect 602 807 636 841
rect 670 807 704 841
rect 738 807 772 841
rect 806 807 840 841
<< locali >>
rect -887 807 -848 841
rect -806 807 -776 841
rect -738 807 -704 841
rect -670 807 -636 841
rect -598 807 -568 841
rect -526 807 -487 841
rect -429 807 -390 841
rect -348 807 -318 841
rect -280 807 -246 841
rect -212 807 -178 841
rect -140 807 -110 841
rect -68 807 -29 841
rect 29 807 68 841
rect 110 807 140 841
rect 178 807 212 841
rect 246 807 280 841
rect 318 807 348 841
rect 390 807 429 841
rect 487 807 526 841
rect 568 807 598 841
rect 636 807 670 841
rect 704 807 738 841
rect 776 807 806 841
rect 848 807 887 841
rect -933 742 -899 773
rect -933 670 -899 700
rect -933 598 -899 632
rect -933 530 -899 564
rect -933 462 -899 492
rect -933 394 -899 420
rect -933 326 -899 348
rect -933 258 -899 276
rect -933 190 -899 204
rect -933 122 -899 132
rect -933 54 -899 60
rect -933 -14 -899 -12
rect -933 -50 -899 -48
rect -933 -122 -899 -116
rect -933 -194 -899 -184
rect -933 -266 -899 -252
rect -933 -338 -899 -320
rect -933 -410 -899 -388
rect -933 -482 -899 -456
rect -933 -554 -899 -524
rect -933 -626 -899 -592
rect -933 -694 -899 -660
rect -933 -762 -899 -732
rect -933 -835 -899 -804
rect -475 742 -441 773
rect -475 670 -441 700
rect -475 598 -441 632
rect -475 530 -441 564
rect -475 462 -441 492
rect -475 394 -441 420
rect -475 326 -441 348
rect -475 258 -441 276
rect -475 190 -441 204
rect -475 122 -441 132
rect -475 54 -441 60
rect -475 -14 -441 -12
rect -475 -50 -441 -48
rect -475 -122 -441 -116
rect -475 -194 -441 -184
rect -475 -266 -441 -252
rect -475 -338 -441 -320
rect -475 -410 -441 -388
rect -475 -482 -441 -456
rect -475 -554 -441 -524
rect -475 -626 -441 -592
rect -475 -694 -441 -660
rect -475 -762 -441 -732
rect -475 -835 -441 -804
rect -17 742 17 773
rect -17 670 17 700
rect -17 598 17 632
rect -17 530 17 564
rect -17 462 17 492
rect -17 394 17 420
rect -17 326 17 348
rect -17 258 17 276
rect -17 190 17 204
rect -17 122 17 132
rect -17 54 17 60
rect -17 -14 17 -12
rect -17 -50 17 -48
rect -17 -122 17 -116
rect -17 -194 17 -184
rect -17 -266 17 -252
rect -17 -338 17 -320
rect -17 -410 17 -388
rect -17 -482 17 -456
rect -17 -554 17 -524
rect -17 -626 17 -592
rect -17 -694 17 -660
rect -17 -762 17 -732
rect -17 -835 17 -804
rect 441 742 475 773
rect 441 670 475 700
rect 441 598 475 632
rect 441 530 475 564
rect 441 462 475 492
rect 441 394 475 420
rect 441 326 475 348
rect 441 258 475 276
rect 441 190 475 204
rect 441 122 475 132
rect 441 54 475 60
rect 441 -14 475 -12
rect 441 -50 475 -48
rect 441 -122 475 -116
rect 441 -194 475 -184
rect 441 -266 475 -252
rect 441 -338 475 -320
rect 441 -410 475 -388
rect 441 -482 475 -456
rect 441 -554 475 -524
rect 441 -626 475 -592
rect 441 -694 475 -660
rect 441 -762 475 -732
rect 441 -835 475 -804
rect 899 742 933 773
rect 899 670 933 700
rect 899 598 933 632
rect 899 530 933 564
rect 899 462 933 492
rect 899 394 933 420
rect 899 326 933 348
rect 899 258 933 276
rect 899 190 933 204
rect 899 122 933 132
rect 899 54 933 60
rect 899 -14 933 -12
rect 899 -50 933 -48
rect 899 -122 933 -116
rect 899 -194 933 -184
rect 899 -266 933 -252
rect 899 -338 933 -320
rect 899 -410 933 -388
rect 899 -482 933 -456
rect 899 -554 933 -524
rect 899 -626 933 -592
rect 899 -694 933 -660
rect 899 -762 933 -732
rect 899 -835 933 -804
<< viali >>
rect -848 807 -840 841
rect -840 807 -814 841
rect -776 807 -772 841
rect -772 807 -742 841
rect -704 807 -670 841
rect -632 807 -602 841
rect -602 807 -598 841
rect -560 807 -534 841
rect -534 807 -526 841
rect -390 807 -382 841
rect -382 807 -356 841
rect -318 807 -314 841
rect -314 807 -284 841
rect -246 807 -212 841
rect -174 807 -144 841
rect -144 807 -140 841
rect -102 807 -76 841
rect -76 807 -68 841
rect 68 807 76 841
rect 76 807 102 841
rect 140 807 144 841
rect 144 807 174 841
rect 212 807 246 841
rect 284 807 314 841
rect 314 807 318 841
rect 356 807 382 841
rect 382 807 390 841
rect 526 807 534 841
rect 534 807 560 841
rect 598 807 602 841
rect 602 807 632 841
rect 670 807 704 841
rect 742 807 772 841
rect 772 807 776 841
rect 814 807 840 841
rect 840 807 848 841
rect -933 734 -899 742
rect -933 708 -899 734
rect -933 666 -899 670
rect -933 636 -899 666
rect -933 564 -899 598
rect -933 496 -899 526
rect -933 492 -899 496
rect -933 428 -899 454
rect -933 420 -899 428
rect -933 360 -899 382
rect -933 348 -899 360
rect -933 292 -899 310
rect -933 276 -899 292
rect -933 224 -899 238
rect -933 204 -899 224
rect -933 156 -899 166
rect -933 132 -899 156
rect -933 88 -899 94
rect -933 60 -899 88
rect -933 20 -899 22
rect -933 -12 -899 20
rect -933 -82 -899 -50
rect -933 -84 -899 -82
rect -933 -150 -899 -122
rect -933 -156 -899 -150
rect -933 -218 -899 -194
rect -933 -228 -899 -218
rect -933 -286 -899 -266
rect -933 -300 -899 -286
rect -933 -354 -899 -338
rect -933 -372 -899 -354
rect -933 -422 -899 -410
rect -933 -444 -899 -422
rect -933 -490 -899 -482
rect -933 -516 -899 -490
rect -933 -558 -899 -554
rect -933 -588 -899 -558
rect -933 -660 -899 -626
rect -933 -728 -899 -698
rect -933 -732 -899 -728
rect -933 -796 -899 -770
rect -933 -804 -899 -796
rect -475 734 -441 742
rect -475 708 -441 734
rect -475 666 -441 670
rect -475 636 -441 666
rect -475 564 -441 598
rect -475 496 -441 526
rect -475 492 -441 496
rect -475 428 -441 454
rect -475 420 -441 428
rect -475 360 -441 382
rect -475 348 -441 360
rect -475 292 -441 310
rect -475 276 -441 292
rect -475 224 -441 238
rect -475 204 -441 224
rect -475 156 -441 166
rect -475 132 -441 156
rect -475 88 -441 94
rect -475 60 -441 88
rect -475 20 -441 22
rect -475 -12 -441 20
rect -475 -82 -441 -50
rect -475 -84 -441 -82
rect -475 -150 -441 -122
rect -475 -156 -441 -150
rect -475 -218 -441 -194
rect -475 -228 -441 -218
rect -475 -286 -441 -266
rect -475 -300 -441 -286
rect -475 -354 -441 -338
rect -475 -372 -441 -354
rect -475 -422 -441 -410
rect -475 -444 -441 -422
rect -475 -490 -441 -482
rect -475 -516 -441 -490
rect -475 -558 -441 -554
rect -475 -588 -441 -558
rect -475 -660 -441 -626
rect -475 -728 -441 -698
rect -475 -732 -441 -728
rect -475 -796 -441 -770
rect -475 -804 -441 -796
rect -17 734 17 742
rect -17 708 17 734
rect -17 666 17 670
rect -17 636 17 666
rect -17 564 17 598
rect -17 496 17 526
rect -17 492 17 496
rect -17 428 17 454
rect -17 420 17 428
rect -17 360 17 382
rect -17 348 17 360
rect -17 292 17 310
rect -17 276 17 292
rect -17 224 17 238
rect -17 204 17 224
rect -17 156 17 166
rect -17 132 17 156
rect -17 88 17 94
rect -17 60 17 88
rect -17 20 17 22
rect -17 -12 17 20
rect -17 -82 17 -50
rect -17 -84 17 -82
rect -17 -150 17 -122
rect -17 -156 17 -150
rect -17 -218 17 -194
rect -17 -228 17 -218
rect -17 -286 17 -266
rect -17 -300 17 -286
rect -17 -354 17 -338
rect -17 -372 17 -354
rect -17 -422 17 -410
rect -17 -444 17 -422
rect -17 -490 17 -482
rect -17 -516 17 -490
rect -17 -558 17 -554
rect -17 -588 17 -558
rect -17 -660 17 -626
rect -17 -728 17 -698
rect -17 -732 17 -728
rect -17 -796 17 -770
rect -17 -804 17 -796
rect 441 734 475 742
rect 441 708 475 734
rect 441 666 475 670
rect 441 636 475 666
rect 441 564 475 598
rect 441 496 475 526
rect 441 492 475 496
rect 441 428 475 454
rect 441 420 475 428
rect 441 360 475 382
rect 441 348 475 360
rect 441 292 475 310
rect 441 276 475 292
rect 441 224 475 238
rect 441 204 475 224
rect 441 156 475 166
rect 441 132 475 156
rect 441 88 475 94
rect 441 60 475 88
rect 441 20 475 22
rect 441 -12 475 20
rect 441 -82 475 -50
rect 441 -84 475 -82
rect 441 -150 475 -122
rect 441 -156 475 -150
rect 441 -218 475 -194
rect 441 -228 475 -218
rect 441 -286 475 -266
rect 441 -300 475 -286
rect 441 -354 475 -338
rect 441 -372 475 -354
rect 441 -422 475 -410
rect 441 -444 475 -422
rect 441 -490 475 -482
rect 441 -516 475 -490
rect 441 -558 475 -554
rect 441 -588 475 -558
rect 441 -660 475 -626
rect 441 -728 475 -698
rect 441 -732 475 -728
rect 441 -796 475 -770
rect 441 -804 475 -796
rect 899 734 933 742
rect 899 708 933 734
rect 899 666 933 670
rect 899 636 933 666
rect 899 564 933 598
rect 899 496 933 526
rect 899 492 933 496
rect 899 428 933 454
rect 899 420 933 428
rect 899 360 933 382
rect 899 348 933 360
rect 899 292 933 310
rect 899 276 933 292
rect 899 224 933 238
rect 899 204 933 224
rect 899 156 933 166
rect 899 132 933 156
rect 899 88 933 94
rect 899 60 933 88
rect 899 20 933 22
rect 899 -12 933 20
rect 899 -82 933 -50
rect 899 -84 933 -82
rect 899 -150 933 -122
rect 899 -156 933 -150
rect 899 -218 933 -194
rect 899 -228 933 -218
rect 899 -286 933 -266
rect 899 -300 933 -286
rect 899 -354 933 -338
rect 899 -372 933 -354
rect 899 -422 933 -410
rect 899 -444 933 -422
rect 899 -490 933 -482
rect 899 -516 933 -490
rect 899 -558 933 -554
rect 899 -588 933 -558
rect 899 -660 933 -626
rect 899 -728 933 -698
rect 899 -732 933 -728
rect 899 -796 933 -770
rect 899 -804 933 -796
<< metal1 >>
rect -883 841 -491 847
rect -883 807 -848 841
rect -814 807 -776 841
rect -742 807 -704 841
rect -670 807 -632 841
rect -598 807 -560 841
rect -526 807 -491 841
rect -883 801 -491 807
rect -425 841 -33 847
rect -425 807 -390 841
rect -356 807 -318 841
rect -284 807 -246 841
rect -212 807 -174 841
rect -140 807 -102 841
rect -68 807 -33 841
rect -425 801 -33 807
rect 33 841 425 847
rect 33 807 68 841
rect 102 807 140 841
rect 174 807 212 841
rect 246 807 284 841
rect 318 807 356 841
rect 390 807 425 841
rect 33 801 425 807
rect 491 841 883 847
rect 491 807 526 841
rect 560 807 598 841
rect 632 807 670 841
rect 704 807 742 841
rect 776 807 814 841
rect 848 807 883 841
rect 491 801 883 807
rect -939 742 -893 769
rect -939 708 -933 742
rect -899 708 -893 742
rect -939 670 -893 708
rect -939 636 -933 670
rect -899 636 -893 670
rect -939 598 -893 636
rect -939 564 -933 598
rect -899 564 -893 598
rect -939 526 -893 564
rect -939 492 -933 526
rect -899 492 -893 526
rect -939 454 -893 492
rect -939 420 -933 454
rect -899 420 -893 454
rect -939 382 -893 420
rect -939 348 -933 382
rect -899 348 -893 382
rect -939 310 -893 348
rect -939 276 -933 310
rect -899 276 -893 310
rect -939 238 -893 276
rect -939 204 -933 238
rect -899 204 -893 238
rect -939 166 -893 204
rect -939 132 -933 166
rect -899 132 -893 166
rect -939 94 -893 132
rect -939 60 -933 94
rect -899 60 -893 94
rect -939 22 -893 60
rect -939 -12 -933 22
rect -899 -12 -893 22
rect -939 -50 -893 -12
rect -939 -84 -933 -50
rect -899 -84 -893 -50
rect -939 -122 -893 -84
rect -939 -156 -933 -122
rect -899 -156 -893 -122
rect -939 -194 -893 -156
rect -939 -228 -933 -194
rect -899 -228 -893 -194
rect -939 -266 -893 -228
rect -939 -300 -933 -266
rect -899 -300 -893 -266
rect -939 -338 -893 -300
rect -939 -372 -933 -338
rect -899 -372 -893 -338
rect -939 -410 -893 -372
rect -939 -444 -933 -410
rect -899 -444 -893 -410
rect -939 -482 -893 -444
rect -939 -516 -933 -482
rect -899 -516 -893 -482
rect -939 -554 -893 -516
rect -939 -588 -933 -554
rect -899 -588 -893 -554
rect -939 -626 -893 -588
rect -939 -660 -933 -626
rect -899 -660 -893 -626
rect -939 -698 -893 -660
rect -939 -732 -933 -698
rect -899 -732 -893 -698
rect -939 -770 -893 -732
rect -939 -804 -933 -770
rect -899 -804 -893 -770
rect -939 -831 -893 -804
rect -481 742 -435 769
rect -481 708 -475 742
rect -441 708 -435 742
rect -481 670 -435 708
rect -481 636 -475 670
rect -441 636 -435 670
rect -481 598 -435 636
rect -481 564 -475 598
rect -441 564 -435 598
rect -481 526 -435 564
rect -481 492 -475 526
rect -441 492 -435 526
rect -481 454 -435 492
rect -481 420 -475 454
rect -441 420 -435 454
rect -481 382 -435 420
rect -481 348 -475 382
rect -441 348 -435 382
rect -481 310 -435 348
rect -481 276 -475 310
rect -441 276 -435 310
rect -481 238 -435 276
rect -481 204 -475 238
rect -441 204 -435 238
rect -481 166 -435 204
rect -481 132 -475 166
rect -441 132 -435 166
rect -481 94 -435 132
rect -481 60 -475 94
rect -441 60 -435 94
rect -481 22 -435 60
rect -481 -12 -475 22
rect -441 -12 -435 22
rect -481 -50 -435 -12
rect -481 -84 -475 -50
rect -441 -84 -435 -50
rect -481 -122 -435 -84
rect -481 -156 -475 -122
rect -441 -156 -435 -122
rect -481 -194 -435 -156
rect -481 -228 -475 -194
rect -441 -228 -435 -194
rect -481 -266 -435 -228
rect -481 -300 -475 -266
rect -441 -300 -435 -266
rect -481 -338 -435 -300
rect -481 -372 -475 -338
rect -441 -372 -435 -338
rect -481 -410 -435 -372
rect -481 -444 -475 -410
rect -441 -444 -435 -410
rect -481 -482 -435 -444
rect -481 -516 -475 -482
rect -441 -516 -435 -482
rect -481 -554 -435 -516
rect -481 -588 -475 -554
rect -441 -588 -435 -554
rect -481 -626 -435 -588
rect -481 -660 -475 -626
rect -441 -660 -435 -626
rect -481 -698 -435 -660
rect -481 -732 -475 -698
rect -441 -732 -435 -698
rect -481 -770 -435 -732
rect -481 -804 -475 -770
rect -441 -804 -435 -770
rect -481 -831 -435 -804
rect -23 742 23 769
rect -23 708 -17 742
rect 17 708 23 742
rect -23 670 23 708
rect -23 636 -17 670
rect 17 636 23 670
rect -23 598 23 636
rect -23 564 -17 598
rect 17 564 23 598
rect -23 526 23 564
rect -23 492 -17 526
rect 17 492 23 526
rect -23 454 23 492
rect -23 420 -17 454
rect 17 420 23 454
rect -23 382 23 420
rect -23 348 -17 382
rect 17 348 23 382
rect -23 310 23 348
rect -23 276 -17 310
rect 17 276 23 310
rect -23 238 23 276
rect -23 204 -17 238
rect 17 204 23 238
rect -23 166 23 204
rect -23 132 -17 166
rect 17 132 23 166
rect -23 94 23 132
rect -23 60 -17 94
rect 17 60 23 94
rect -23 22 23 60
rect -23 -12 -17 22
rect 17 -12 23 22
rect -23 -50 23 -12
rect -23 -84 -17 -50
rect 17 -84 23 -50
rect -23 -122 23 -84
rect -23 -156 -17 -122
rect 17 -156 23 -122
rect -23 -194 23 -156
rect -23 -228 -17 -194
rect 17 -228 23 -194
rect -23 -266 23 -228
rect -23 -300 -17 -266
rect 17 -300 23 -266
rect -23 -338 23 -300
rect -23 -372 -17 -338
rect 17 -372 23 -338
rect -23 -410 23 -372
rect -23 -444 -17 -410
rect 17 -444 23 -410
rect -23 -482 23 -444
rect -23 -516 -17 -482
rect 17 -516 23 -482
rect -23 -554 23 -516
rect -23 -588 -17 -554
rect 17 -588 23 -554
rect -23 -626 23 -588
rect -23 -660 -17 -626
rect 17 -660 23 -626
rect -23 -698 23 -660
rect -23 -732 -17 -698
rect 17 -732 23 -698
rect -23 -770 23 -732
rect -23 -804 -17 -770
rect 17 -804 23 -770
rect -23 -831 23 -804
rect 435 742 481 769
rect 435 708 441 742
rect 475 708 481 742
rect 435 670 481 708
rect 435 636 441 670
rect 475 636 481 670
rect 435 598 481 636
rect 435 564 441 598
rect 475 564 481 598
rect 435 526 481 564
rect 435 492 441 526
rect 475 492 481 526
rect 435 454 481 492
rect 435 420 441 454
rect 475 420 481 454
rect 435 382 481 420
rect 435 348 441 382
rect 475 348 481 382
rect 435 310 481 348
rect 435 276 441 310
rect 475 276 481 310
rect 435 238 481 276
rect 435 204 441 238
rect 475 204 481 238
rect 435 166 481 204
rect 435 132 441 166
rect 475 132 481 166
rect 435 94 481 132
rect 435 60 441 94
rect 475 60 481 94
rect 435 22 481 60
rect 435 -12 441 22
rect 475 -12 481 22
rect 435 -50 481 -12
rect 435 -84 441 -50
rect 475 -84 481 -50
rect 435 -122 481 -84
rect 435 -156 441 -122
rect 475 -156 481 -122
rect 435 -194 481 -156
rect 435 -228 441 -194
rect 475 -228 481 -194
rect 435 -266 481 -228
rect 435 -300 441 -266
rect 475 -300 481 -266
rect 435 -338 481 -300
rect 435 -372 441 -338
rect 475 -372 481 -338
rect 435 -410 481 -372
rect 435 -444 441 -410
rect 475 -444 481 -410
rect 435 -482 481 -444
rect 435 -516 441 -482
rect 475 -516 481 -482
rect 435 -554 481 -516
rect 435 -588 441 -554
rect 475 -588 481 -554
rect 435 -626 481 -588
rect 435 -660 441 -626
rect 475 -660 481 -626
rect 435 -698 481 -660
rect 435 -732 441 -698
rect 475 -732 481 -698
rect 435 -770 481 -732
rect 435 -804 441 -770
rect 475 -804 481 -770
rect 435 -831 481 -804
rect 893 742 939 769
rect 893 708 899 742
rect 933 708 939 742
rect 893 670 939 708
rect 893 636 899 670
rect 933 636 939 670
rect 893 598 939 636
rect 893 564 899 598
rect 933 564 939 598
rect 893 526 939 564
rect 893 492 899 526
rect 933 492 939 526
rect 893 454 939 492
rect 893 420 899 454
rect 933 420 939 454
rect 893 382 939 420
rect 893 348 899 382
rect 933 348 939 382
rect 893 310 939 348
rect 893 276 899 310
rect 933 276 939 310
rect 893 238 939 276
rect 893 204 899 238
rect 933 204 939 238
rect 893 166 939 204
rect 893 132 899 166
rect 933 132 939 166
rect 893 94 939 132
rect 893 60 899 94
rect 933 60 939 94
rect 893 22 939 60
rect 893 -12 899 22
rect 933 -12 939 22
rect 893 -50 939 -12
rect 893 -84 899 -50
rect 933 -84 939 -50
rect 893 -122 939 -84
rect 893 -156 899 -122
rect 933 -156 939 -122
rect 893 -194 939 -156
rect 893 -228 899 -194
rect 933 -228 939 -194
rect 893 -266 939 -228
rect 893 -300 899 -266
rect 933 -300 939 -266
rect 893 -338 939 -300
rect 893 -372 899 -338
rect 933 -372 939 -338
rect 893 -410 939 -372
rect 893 -444 899 -410
rect 933 -444 939 -410
rect 893 -482 939 -444
rect 893 -516 899 -482
rect 933 -516 939 -482
rect 893 -554 939 -516
rect 893 -588 899 -554
rect 933 -588 939 -554
rect 893 -626 939 -588
rect 893 -660 899 -626
rect 933 -660 939 -626
rect 893 -698 939 -660
rect 893 -732 899 -698
rect 933 -732 939 -698
rect 893 -770 939 -732
rect 893 -804 899 -770
rect 933 -804 939 -770
rect 893 -831 939 -804
<< end >>
