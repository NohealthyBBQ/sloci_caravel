magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal4 >>
rect -951 438 951 500
rect -951 202 695 438
rect 931 202 951 438
rect -951 118 951 202
rect -951 -118 695 118
rect 931 -118 951 118
rect -951 -202 951 -118
rect -951 -438 695 -202
rect 931 -438 951 -202
rect -951 -500 951 -438
<< via4 >>
rect 695 202 931 438
rect 695 -118 931 118
rect 695 -438 931 -202
<< mimcap2 >>
rect -851 278 349 400
rect -851 -278 -689 278
rect 187 -278 349 278
rect -851 -400 349 -278
<< mimcap2contact >>
rect -689 -278 187 278
<< metal5 >>
rect 653 438 973 501
rect -835 278 333 384
rect -835 -278 -689 278
rect 187 -278 333 278
rect -835 -384 333 -278
rect 653 202 695 438
rect 931 202 973 438
rect 653 118 973 202
rect 653 -118 695 118
rect 931 -118 973 118
rect 653 -202 973 -118
rect 653 -438 695 -202
rect 931 -438 973 -202
rect 653 -501 973 -438
<< properties >>
string FIXED_BBOX -951 -500 449 500
<< end >>
