magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -297 4741 297 4827
rect -297 -4741 -211 4741
rect 211 -4741 297 4741
rect -297 -4827 297 -4741
<< psubdiff >>
rect -271 4767 -153 4801
rect -119 4767 -85 4801
rect -51 4767 -17 4801
rect 17 4767 51 4801
rect 85 4767 119 4801
rect 153 4767 271 4801
rect -271 4675 -237 4767
rect 237 4675 271 4767
rect -271 4607 -237 4641
rect -271 4539 -237 4573
rect -271 4471 -237 4505
rect -271 4403 -237 4437
rect -271 4335 -237 4369
rect -271 4267 -237 4301
rect -271 4199 -237 4233
rect -271 4131 -237 4165
rect -271 4063 -237 4097
rect -271 3995 -237 4029
rect -271 3927 -237 3961
rect -271 3859 -237 3893
rect -271 3791 -237 3825
rect -271 3723 -237 3757
rect -271 3655 -237 3689
rect -271 3587 -237 3621
rect -271 3519 -237 3553
rect -271 3451 -237 3485
rect -271 3383 -237 3417
rect -271 3315 -237 3349
rect -271 3247 -237 3281
rect -271 3179 -237 3213
rect -271 3111 -237 3145
rect -271 3043 -237 3077
rect -271 2975 -237 3009
rect -271 2907 -237 2941
rect -271 2839 -237 2873
rect -271 2771 -237 2805
rect -271 2703 -237 2737
rect -271 2635 -237 2669
rect -271 2567 -237 2601
rect -271 2499 -237 2533
rect -271 2431 -237 2465
rect -271 2363 -237 2397
rect -271 2295 -237 2329
rect -271 2227 -237 2261
rect -271 2159 -237 2193
rect -271 2091 -237 2125
rect -271 2023 -237 2057
rect -271 1955 -237 1989
rect -271 1887 -237 1921
rect -271 1819 -237 1853
rect -271 1751 -237 1785
rect -271 1683 -237 1717
rect -271 1615 -237 1649
rect -271 1547 -237 1581
rect -271 1479 -237 1513
rect -271 1411 -237 1445
rect -271 1343 -237 1377
rect -271 1275 -237 1309
rect -271 1207 -237 1241
rect -271 1139 -237 1173
rect -271 1071 -237 1105
rect -271 1003 -237 1037
rect -271 935 -237 969
rect -271 867 -237 901
rect -271 799 -237 833
rect -271 731 -237 765
rect -271 663 -237 697
rect -271 595 -237 629
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect -271 -629 -237 -595
rect -271 -697 -237 -663
rect -271 -765 -237 -731
rect -271 -833 -237 -799
rect -271 -901 -237 -867
rect -271 -969 -237 -935
rect -271 -1037 -237 -1003
rect -271 -1105 -237 -1071
rect -271 -1173 -237 -1139
rect -271 -1241 -237 -1207
rect -271 -1309 -237 -1275
rect -271 -1377 -237 -1343
rect -271 -1445 -237 -1411
rect -271 -1513 -237 -1479
rect -271 -1581 -237 -1547
rect -271 -1649 -237 -1615
rect -271 -1717 -237 -1683
rect -271 -1785 -237 -1751
rect -271 -1853 -237 -1819
rect -271 -1921 -237 -1887
rect -271 -1989 -237 -1955
rect -271 -2057 -237 -2023
rect -271 -2125 -237 -2091
rect -271 -2193 -237 -2159
rect -271 -2261 -237 -2227
rect -271 -2329 -237 -2295
rect -271 -2397 -237 -2363
rect -271 -2465 -237 -2431
rect -271 -2533 -237 -2499
rect -271 -2601 -237 -2567
rect -271 -2669 -237 -2635
rect -271 -2737 -237 -2703
rect -271 -2805 -237 -2771
rect -271 -2873 -237 -2839
rect -271 -2941 -237 -2907
rect -271 -3009 -237 -2975
rect -271 -3077 -237 -3043
rect -271 -3145 -237 -3111
rect -271 -3213 -237 -3179
rect -271 -3281 -237 -3247
rect -271 -3349 -237 -3315
rect -271 -3417 -237 -3383
rect -271 -3485 -237 -3451
rect -271 -3553 -237 -3519
rect -271 -3621 -237 -3587
rect -271 -3689 -237 -3655
rect -271 -3757 -237 -3723
rect -271 -3825 -237 -3791
rect -271 -3893 -237 -3859
rect -271 -3961 -237 -3927
rect -271 -4029 -237 -3995
rect -271 -4097 -237 -4063
rect -271 -4165 -237 -4131
rect -271 -4233 -237 -4199
rect -271 -4301 -237 -4267
rect -271 -4369 -237 -4335
rect -271 -4437 -237 -4403
rect -271 -4505 -237 -4471
rect -271 -4573 -237 -4539
rect -271 -4641 -237 -4607
rect 237 4607 271 4641
rect 237 4539 271 4573
rect 237 4471 271 4505
rect 237 4403 271 4437
rect 237 4335 271 4369
rect 237 4267 271 4301
rect 237 4199 271 4233
rect 237 4131 271 4165
rect 237 4063 271 4097
rect 237 3995 271 4029
rect 237 3927 271 3961
rect 237 3859 271 3893
rect 237 3791 271 3825
rect 237 3723 271 3757
rect 237 3655 271 3689
rect 237 3587 271 3621
rect 237 3519 271 3553
rect 237 3451 271 3485
rect 237 3383 271 3417
rect 237 3315 271 3349
rect 237 3247 271 3281
rect 237 3179 271 3213
rect 237 3111 271 3145
rect 237 3043 271 3077
rect 237 2975 271 3009
rect 237 2907 271 2941
rect 237 2839 271 2873
rect 237 2771 271 2805
rect 237 2703 271 2737
rect 237 2635 271 2669
rect 237 2567 271 2601
rect 237 2499 271 2533
rect 237 2431 271 2465
rect 237 2363 271 2397
rect 237 2295 271 2329
rect 237 2227 271 2261
rect 237 2159 271 2193
rect 237 2091 271 2125
rect 237 2023 271 2057
rect 237 1955 271 1989
rect 237 1887 271 1921
rect 237 1819 271 1853
rect 237 1751 271 1785
rect 237 1683 271 1717
rect 237 1615 271 1649
rect 237 1547 271 1581
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1207 271 1241
rect 237 1139 271 1173
rect 237 1071 271 1105
rect 237 1003 271 1037
rect 237 935 271 969
rect 237 867 271 901
rect 237 799 271 833
rect 237 731 271 765
rect 237 663 271 697
rect 237 595 271 629
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect 237 -629 271 -595
rect 237 -697 271 -663
rect 237 -765 271 -731
rect 237 -833 271 -799
rect 237 -901 271 -867
rect 237 -969 271 -935
rect 237 -1037 271 -1003
rect 237 -1105 271 -1071
rect 237 -1173 271 -1139
rect 237 -1241 271 -1207
rect 237 -1309 271 -1275
rect 237 -1377 271 -1343
rect 237 -1445 271 -1411
rect 237 -1513 271 -1479
rect 237 -1581 271 -1547
rect 237 -1649 271 -1615
rect 237 -1717 271 -1683
rect 237 -1785 271 -1751
rect 237 -1853 271 -1819
rect 237 -1921 271 -1887
rect 237 -1989 271 -1955
rect 237 -2057 271 -2023
rect 237 -2125 271 -2091
rect 237 -2193 271 -2159
rect 237 -2261 271 -2227
rect 237 -2329 271 -2295
rect 237 -2397 271 -2363
rect 237 -2465 271 -2431
rect 237 -2533 271 -2499
rect 237 -2601 271 -2567
rect 237 -2669 271 -2635
rect 237 -2737 271 -2703
rect 237 -2805 271 -2771
rect 237 -2873 271 -2839
rect 237 -2941 271 -2907
rect 237 -3009 271 -2975
rect 237 -3077 271 -3043
rect 237 -3145 271 -3111
rect 237 -3213 271 -3179
rect 237 -3281 271 -3247
rect 237 -3349 271 -3315
rect 237 -3417 271 -3383
rect 237 -3485 271 -3451
rect 237 -3553 271 -3519
rect 237 -3621 271 -3587
rect 237 -3689 271 -3655
rect 237 -3757 271 -3723
rect 237 -3825 271 -3791
rect 237 -3893 271 -3859
rect 237 -3961 271 -3927
rect 237 -4029 271 -3995
rect 237 -4097 271 -4063
rect 237 -4165 271 -4131
rect 237 -4233 271 -4199
rect 237 -4301 271 -4267
rect 237 -4369 271 -4335
rect 237 -4437 271 -4403
rect 237 -4505 271 -4471
rect 237 -4573 271 -4539
rect 237 -4641 271 -4607
rect -271 -4767 -237 -4675
rect 237 -4767 271 -4675
rect -271 -4801 -153 -4767
rect -119 -4801 -85 -4767
rect -51 -4801 -17 -4767
rect 17 -4801 51 -4767
rect 85 -4801 119 -4767
rect 153 -4801 271 -4767
<< psubdiffcont >>
rect -153 4767 -119 4801
rect -85 4767 -51 4801
rect -17 4767 17 4801
rect 51 4767 85 4801
rect 119 4767 153 4801
rect -271 4641 -237 4675
rect -271 4573 -237 4607
rect -271 4505 -237 4539
rect -271 4437 -237 4471
rect -271 4369 -237 4403
rect -271 4301 -237 4335
rect -271 4233 -237 4267
rect -271 4165 -237 4199
rect -271 4097 -237 4131
rect -271 4029 -237 4063
rect -271 3961 -237 3995
rect -271 3893 -237 3927
rect -271 3825 -237 3859
rect -271 3757 -237 3791
rect -271 3689 -237 3723
rect -271 3621 -237 3655
rect -271 3553 -237 3587
rect -271 3485 -237 3519
rect -271 3417 -237 3451
rect -271 3349 -237 3383
rect -271 3281 -237 3315
rect -271 3213 -237 3247
rect -271 3145 -237 3179
rect -271 3077 -237 3111
rect -271 3009 -237 3043
rect -271 2941 -237 2975
rect -271 2873 -237 2907
rect -271 2805 -237 2839
rect -271 2737 -237 2771
rect -271 2669 -237 2703
rect -271 2601 -237 2635
rect -271 2533 -237 2567
rect -271 2465 -237 2499
rect -271 2397 -237 2431
rect -271 2329 -237 2363
rect -271 2261 -237 2295
rect -271 2193 -237 2227
rect -271 2125 -237 2159
rect -271 2057 -237 2091
rect -271 1989 -237 2023
rect -271 1921 -237 1955
rect -271 1853 -237 1887
rect -271 1785 -237 1819
rect -271 1717 -237 1751
rect -271 1649 -237 1683
rect -271 1581 -237 1615
rect -271 1513 -237 1547
rect -271 1445 -237 1479
rect -271 1377 -237 1411
rect -271 1309 -237 1343
rect -271 1241 -237 1275
rect -271 1173 -237 1207
rect -271 1105 -237 1139
rect -271 1037 -237 1071
rect -271 969 -237 1003
rect -271 901 -237 935
rect -271 833 -237 867
rect -271 765 -237 799
rect -271 697 -237 731
rect -271 629 -237 663
rect -271 561 -237 595
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect -271 -595 -237 -561
rect -271 -663 -237 -629
rect -271 -731 -237 -697
rect -271 -799 -237 -765
rect -271 -867 -237 -833
rect -271 -935 -237 -901
rect -271 -1003 -237 -969
rect -271 -1071 -237 -1037
rect -271 -1139 -237 -1105
rect -271 -1207 -237 -1173
rect -271 -1275 -237 -1241
rect -271 -1343 -237 -1309
rect -271 -1411 -237 -1377
rect -271 -1479 -237 -1445
rect -271 -1547 -237 -1513
rect -271 -1615 -237 -1581
rect -271 -1683 -237 -1649
rect -271 -1751 -237 -1717
rect -271 -1819 -237 -1785
rect -271 -1887 -237 -1853
rect -271 -1955 -237 -1921
rect -271 -2023 -237 -1989
rect -271 -2091 -237 -2057
rect -271 -2159 -237 -2125
rect -271 -2227 -237 -2193
rect -271 -2295 -237 -2261
rect -271 -2363 -237 -2329
rect -271 -2431 -237 -2397
rect -271 -2499 -237 -2465
rect -271 -2567 -237 -2533
rect -271 -2635 -237 -2601
rect -271 -2703 -237 -2669
rect -271 -2771 -237 -2737
rect -271 -2839 -237 -2805
rect -271 -2907 -237 -2873
rect -271 -2975 -237 -2941
rect -271 -3043 -237 -3009
rect -271 -3111 -237 -3077
rect -271 -3179 -237 -3145
rect -271 -3247 -237 -3213
rect -271 -3315 -237 -3281
rect -271 -3383 -237 -3349
rect -271 -3451 -237 -3417
rect -271 -3519 -237 -3485
rect -271 -3587 -237 -3553
rect -271 -3655 -237 -3621
rect -271 -3723 -237 -3689
rect -271 -3791 -237 -3757
rect -271 -3859 -237 -3825
rect -271 -3927 -237 -3893
rect -271 -3995 -237 -3961
rect -271 -4063 -237 -4029
rect -271 -4131 -237 -4097
rect -271 -4199 -237 -4165
rect -271 -4267 -237 -4233
rect -271 -4335 -237 -4301
rect -271 -4403 -237 -4369
rect -271 -4471 -237 -4437
rect -271 -4539 -237 -4505
rect -271 -4607 -237 -4573
rect -271 -4675 -237 -4641
rect 237 4641 271 4675
rect 237 4573 271 4607
rect 237 4505 271 4539
rect 237 4437 271 4471
rect 237 4369 271 4403
rect 237 4301 271 4335
rect 237 4233 271 4267
rect 237 4165 271 4199
rect 237 4097 271 4131
rect 237 4029 271 4063
rect 237 3961 271 3995
rect 237 3893 271 3927
rect 237 3825 271 3859
rect 237 3757 271 3791
rect 237 3689 271 3723
rect 237 3621 271 3655
rect 237 3553 271 3587
rect 237 3485 271 3519
rect 237 3417 271 3451
rect 237 3349 271 3383
rect 237 3281 271 3315
rect 237 3213 271 3247
rect 237 3145 271 3179
rect 237 3077 271 3111
rect 237 3009 271 3043
rect 237 2941 271 2975
rect 237 2873 271 2907
rect 237 2805 271 2839
rect 237 2737 271 2771
rect 237 2669 271 2703
rect 237 2601 271 2635
rect 237 2533 271 2567
rect 237 2465 271 2499
rect 237 2397 271 2431
rect 237 2329 271 2363
rect 237 2261 271 2295
rect 237 2193 271 2227
rect 237 2125 271 2159
rect 237 2057 271 2091
rect 237 1989 271 2023
rect 237 1921 271 1955
rect 237 1853 271 1887
rect 237 1785 271 1819
rect 237 1717 271 1751
rect 237 1649 271 1683
rect 237 1581 271 1615
rect 237 1513 271 1547
rect 237 1445 271 1479
rect 237 1377 271 1411
rect 237 1309 271 1343
rect 237 1241 271 1275
rect 237 1173 271 1207
rect 237 1105 271 1139
rect 237 1037 271 1071
rect 237 969 271 1003
rect 237 901 271 935
rect 237 833 271 867
rect 237 765 271 799
rect 237 697 271 731
rect 237 629 271 663
rect 237 561 271 595
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect 237 -595 271 -561
rect 237 -663 271 -629
rect 237 -731 271 -697
rect 237 -799 271 -765
rect 237 -867 271 -833
rect 237 -935 271 -901
rect 237 -1003 271 -969
rect 237 -1071 271 -1037
rect 237 -1139 271 -1105
rect 237 -1207 271 -1173
rect 237 -1275 271 -1241
rect 237 -1343 271 -1309
rect 237 -1411 271 -1377
rect 237 -1479 271 -1445
rect 237 -1547 271 -1513
rect 237 -1615 271 -1581
rect 237 -1683 271 -1649
rect 237 -1751 271 -1717
rect 237 -1819 271 -1785
rect 237 -1887 271 -1853
rect 237 -1955 271 -1921
rect 237 -2023 271 -1989
rect 237 -2091 271 -2057
rect 237 -2159 271 -2125
rect 237 -2227 271 -2193
rect 237 -2295 271 -2261
rect 237 -2363 271 -2329
rect 237 -2431 271 -2397
rect 237 -2499 271 -2465
rect 237 -2567 271 -2533
rect 237 -2635 271 -2601
rect 237 -2703 271 -2669
rect 237 -2771 271 -2737
rect 237 -2839 271 -2805
rect 237 -2907 271 -2873
rect 237 -2975 271 -2941
rect 237 -3043 271 -3009
rect 237 -3111 271 -3077
rect 237 -3179 271 -3145
rect 237 -3247 271 -3213
rect 237 -3315 271 -3281
rect 237 -3383 271 -3349
rect 237 -3451 271 -3417
rect 237 -3519 271 -3485
rect 237 -3587 271 -3553
rect 237 -3655 271 -3621
rect 237 -3723 271 -3689
rect 237 -3791 271 -3757
rect 237 -3859 271 -3825
rect 237 -3927 271 -3893
rect 237 -3995 271 -3961
rect 237 -4063 271 -4029
rect 237 -4131 271 -4097
rect 237 -4199 271 -4165
rect 237 -4267 271 -4233
rect 237 -4335 271 -4301
rect 237 -4403 271 -4369
rect 237 -4471 271 -4437
rect 237 -4539 271 -4505
rect 237 -4607 271 -4573
rect 237 -4675 271 -4641
rect -153 -4801 -119 -4767
rect -85 -4801 -51 -4767
rect -17 -4801 17 -4767
rect 51 -4801 85 -4767
rect 119 -4801 153 -4767
<< xpolycontact >>
rect -141 4239 141 4671
rect -141 -4671 141 -4239
<< ppolyres >>
rect -141 -4239 141 4239
<< locali >>
rect -271 4767 -153 4801
rect -119 4767 -85 4801
rect -51 4767 -17 4801
rect 17 4767 51 4801
rect 85 4767 119 4801
rect 153 4767 271 4801
rect -271 4675 -237 4767
rect 237 4675 271 4767
rect -271 4607 -237 4641
rect -271 4539 -237 4573
rect -271 4471 -237 4505
rect -271 4403 -237 4437
rect -271 4335 -237 4369
rect -271 4267 -237 4301
rect 237 4607 271 4641
rect 237 4539 271 4573
rect 237 4471 271 4505
rect 237 4403 271 4437
rect 237 4335 271 4369
rect 237 4267 271 4301
rect -271 4199 -237 4233
rect -271 4131 -237 4165
rect -271 4063 -237 4097
rect -271 3995 -237 4029
rect -271 3927 -237 3961
rect -271 3859 -237 3893
rect -271 3791 -237 3825
rect -271 3723 -237 3757
rect -271 3655 -237 3689
rect -271 3587 -237 3621
rect -271 3519 -237 3553
rect -271 3451 -237 3485
rect -271 3383 -237 3417
rect -271 3315 -237 3349
rect -271 3247 -237 3281
rect -271 3179 -237 3213
rect -271 3111 -237 3145
rect -271 3043 -237 3077
rect -271 2975 -237 3009
rect -271 2907 -237 2941
rect -271 2839 -237 2873
rect -271 2771 -237 2805
rect -271 2703 -237 2737
rect -271 2635 -237 2669
rect -271 2567 -237 2601
rect -271 2499 -237 2533
rect -271 2431 -237 2465
rect -271 2363 -237 2397
rect -271 2295 -237 2329
rect -271 2227 -237 2261
rect -271 2159 -237 2193
rect -271 2091 -237 2125
rect -271 2023 -237 2057
rect -271 1955 -237 1989
rect -271 1887 -237 1921
rect -271 1819 -237 1853
rect -271 1751 -237 1785
rect -271 1683 -237 1717
rect -271 1615 -237 1649
rect -271 1547 -237 1581
rect -271 1479 -237 1513
rect -271 1411 -237 1445
rect -271 1343 -237 1377
rect -271 1275 -237 1309
rect -271 1207 -237 1241
rect -271 1139 -237 1173
rect -271 1071 -237 1105
rect -271 1003 -237 1037
rect -271 935 -237 969
rect -271 867 -237 901
rect -271 799 -237 833
rect -271 731 -237 765
rect -271 663 -237 697
rect -271 595 -237 629
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect -271 -629 -237 -595
rect -271 -697 -237 -663
rect -271 -765 -237 -731
rect -271 -833 -237 -799
rect -271 -901 -237 -867
rect -271 -969 -237 -935
rect -271 -1037 -237 -1003
rect -271 -1105 -237 -1071
rect -271 -1173 -237 -1139
rect -271 -1241 -237 -1207
rect -271 -1309 -237 -1275
rect -271 -1377 -237 -1343
rect -271 -1445 -237 -1411
rect -271 -1513 -237 -1479
rect -271 -1581 -237 -1547
rect -271 -1649 -237 -1615
rect -271 -1717 -237 -1683
rect -271 -1785 -237 -1751
rect -271 -1853 -237 -1819
rect -271 -1921 -237 -1887
rect -271 -1989 -237 -1955
rect -271 -2057 -237 -2023
rect -271 -2125 -237 -2091
rect -271 -2193 -237 -2159
rect -271 -2261 -237 -2227
rect -271 -2329 -237 -2295
rect -271 -2397 -237 -2363
rect -271 -2465 -237 -2431
rect -271 -2533 -237 -2499
rect -271 -2601 -237 -2567
rect -271 -2669 -237 -2635
rect -271 -2737 -237 -2703
rect -271 -2805 -237 -2771
rect -271 -2873 -237 -2839
rect -271 -2941 -237 -2907
rect -271 -3009 -237 -2975
rect -271 -3077 -237 -3043
rect -271 -3145 -237 -3111
rect -271 -3213 -237 -3179
rect -271 -3281 -237 -3247
rect -271 -3349 -237 -3315
rect -271 -3417 -237 -3383
rect -271 -3485 -237 -3451
rect -271 -3553 -237 -3519
rect -271 -3621 -237 -3587
rect -271 -3689 -237 -3655
rect -271 -3757 -237 -3723
rect -271 -3825 -237 -3791
rect -271 -3893 -237 -3859
rect -271 -3961 -237 -3927
rect -271 -4029 -237 -3995
rect -271 -4097 -237 -4063
rect -271 -4165 -237 -4131
rect -271 -4233 -237 -4199
rect 237 4199 271 4233
rect 237 4131 271 4165
rect 237 4063 271 4097
rect 237 3995 271 4029
rect 237 3927 271 3961
rect 237 3859 271 3893
rect 237 3791 271 3825
rect 237 3723 271 3757
rect 237 3655 271 3689
rect 237 3587 271 3621
rect 237 3519 271 3553
rect 237 3451 271 3485
rect 237 3383 271 3417
rect 237 3315 271 3349
rect 237 3247 271 3281
rect 237 3179 271 3213
rect 237 3111 271 3145
rect 237 3043 271 3077
rect 237 2975 271 3009
rect 237 2907 271 2941
rect 237 2839 271 2873
rect 237 2771 271 2805
rect 237 2703 271 2737
rect 237 2635 271 2669
rect 237 2567 271 2601
rect 237 2499 271 2533
rect 237 2431 271 2465
rect 237 2363 271 2397
rect 237 2295 271 2329
rect 237 2227 271 2261
rect 237 2159 271 2193
rect 237 2091 271 2125
rect 237 2023 271 2057
rect 237 1955 271 1989
rect 237 1887 271 1921
rect 237 1819 271 1853
rect 237 1751 271 1785
rect 237 1683 271 1717
rect 237 1615 271 1649
rect 237 1547 271 1581
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1207 271 1241
rect 237 1139 271 1173
rect 237 1071 271 1105
rect 237 1003 271 1037
rect 237 935 271 969
rect 237 867 271 901
rect 237 799 271 833
rect 237 731 271 765
rect 237 663 271 697
rect 237 595 271 629
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect 237 -629 271 -595
rect 237 -697 271 -663
rect 237 -765 271 -731
rect 237 -833 271 -799
rect 237 -901 271 -867
rect 237 -969 271 -935
rect 237 -1037 271 -1003
rect 237 -1105 271 -1071
rect 237 -1173 271 -1139
rect 237 -1241 271 -1207
rect 237 -1309 271 -1275
rect 237 -1377 271 -1343
rect 237 -1445 271 -1411
rect 237 -1513 271 -1479
rect 237 -1581 271 -1547
rect 237 -1649 271 -1615
rect 237 -1717 271 -1683
rect 237 -1785 271 -1751
rect 237 -1853 271 -1819
rect 237 -1921 271 -1887
rect 237 -1989 271 -1955
rect 237 -2057 271 -2023
rect 237 -2125 271 -2091
rect 237 -2193 271 -2159
rect 237 -2261 271 -2227
rect 237 -2329 271 -2295
rect 237 -2397 271 -2363
rect 237 -2465 271 -2431
rect 237 -2533 271 -2499
rect 237 -2601 271 -2567
rect 237 -2669 271 -2635
rect 237 -2737 271 -2703
rect 237 -2805 271 -2771
rect 237 -2873 271 -2839
rect 237 -2941 271 -2907
rect 237 -3009 271 -2975
rect 237 -3077 271 -3043
rect 237 -3145 271 -3111
rect 237 -3213 271 -3179
rect 237 -3281 271 -3247
rect 237 -3349 271 -3315
rect 237 -3417 271 -3383
rect 237 -3485 271 -3451
rect 237 -3553 271 -3519
rect 237 -3621 271 -3587
rect 237 -3689 271 -3655
rect 237 -3757 271 -3723
rect 237 -3825 271 -3791
rect 237 -3893 271 -3859
rect 237 -3961 271 -3927
rect 237 -4029 271 -3995
rect 237 -4097 271 -4063
rect 237 -4165 271 -4131
rect 237 -4233 271 -4199
rect -271 -4301 -237 -4267
rect -271 -4369 -237 -4335
rect -271 -4437 -237 -4403
rect -271 -4505 -237 -4471
rect -271 -4573 -237 -4539
rect -271 -4641 -237 -4607
rect 237 -4301 271 -4267
rect 237 -4369 271 -4335
rect 237 -4437 271 -4403
rect 237 -4505 271 -4471
rect 237 -4573 271 -4539
rect 237 -4641 271 -4607
rect -271 -4767 -237 -4675
rect 237 -4767 271 -4675
rect -271 -4801 -153 -4767
rect -119 -4801 -85 -4767
rect -51 -4801 -17 -4767
rect 17 -4801 51 -4767
rect 85 -4801 119 -4767
rect 153 -4801 271 -4767
<< viali >>
rect -125 4257 125 4651
rect -125 -4652 125 -4258
<< metal1 >>
rect -131 4651 131 4665
rect -131 4257 -125 4651
rect 125 4257 131 4651
rect -131 4244 131 4257
rect -131 -4258 131 -4244
rect -131 -4652 -125 -4258
rect 125 -4652 131 -4258
rect -131 -4665 131 -4652
<< properties >>
string FIXED_BBOX -254 -4784 254 4784
<< end >>
