magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -441 1262 441 1348
rect -441 -1262 -355 1262
rect 355 -1262 441 1262
rect -441 -1348 441 -1262
<< psubdiff >>
rect -415 1288 -289 1322
rect -255 1288 -221 1322
rect -187 1288 -153 1322
rect -119 1288 -85 1322
rect -51 1288 -17 1322
rect 17 1288 51 1322
rect 85 1288 119 1322
rect 153 1288 187 1322
rect 221 1288 255 1322
rect 289 1288 415 1322
rect -415 1207 -381 1288
rect 381 1207 415 1288
rect -415 1139 -381 1173
rect -415 1071 -381 1105
rect -415 1003 -381 1037
rect -415 935 -381 969
rect -415 867 -381 901
rect -415 799 -381 833
rect -415 731 -381 765
rect -415 663 -381 697
rect -415 595 -381 629
rect -415 527 -381 561
rect -415 459 -381 493
rect -415 391 -381 425
rect -415 323 -381 357
rect -415 255 -381 289
rect -415 187 -381 221
rect -415 119 -381 153
rect -415 51 -381 85
rect -415 -17 -381 17
rect -415 -85 -381 -51
rect -415 -153 -381 -119
rect -415 -221 -381 -187
rect -415 -289 -381 -255
rect -415 -357 -381 -323
rect -415 -425 -381 -391
rect -415 -493 -381 -459
rect -415 -561 -381 -527
rect -415 -629 -381 -595
rect -415 -697 -381 -663
rect -415 -765 -381 -731
rect -415 -833 -381 -799
rect -415 -901 -381 -867
rect -415 -969 -381 -935
rect -415 -1037 -381 -1003
rect -415 -1105 -381 -1071
rect -415 -1173 -381 -1139
rect 381 1139 415 1173
rect 381 1071 415 1105
rect 381 1003 415 1037
rect 381 935 415 969
rect 381 867 415 901
rect 381 799 415 833
rect 381 731 415 765
rect 381 663 415 697
rect 381 595 415 629
rect 381 527 415 561
rect 381 459 415 493
rect 381 391 415 425
rect 381 323 415 357
rect 381 255 415 289
rect 381 187 415 221
rect 381 119 415 153
rect 381 51 415 85
rect 381 -17 415 17
rect 381 -85 415 -51
rect 381 -153 415 -119
rect 381 -221 415 -187
rect 381 -289 415 -255
rect 381 -357 415 -323
rect 381 -425 415 -391
rect 381 -493 415 -459
rect 381 -561 415 -527
rect 381 -629 415 -595
rect 381 -697 415 -663
rect 381 -765 415 -731
rect 381 -833 415 -799
rect 381 -901 415 -867
rect 381 -969 415 -935
rect 381 -1037 415 -1003
rect 381 -1105 415 -1071
rect 381 -1173 415 -1139
rect -415 -1288 -381 -1207
rect 381 -1288 415 -1207
rect -415 -1322 -289 -1288
rect -255 -1322 -221 -1288
rect -187 -1322 -153 -1288
rect -119 -1322 -85 -1288
rect -51 -1322 -17 -1288
rect 17 -1322 51 -1288
rect 85 -1322 119 -1288
rect 153 -1322 187 -1288
rect 221 -1322 255 -1288
rect 289 -1322 415 -1288
<< psubdiffcont >>
rect -289 1288 -255 1322
rect -221 1288 -187 1322
rect -153 1288 -119 1322
rect -85 1288 -51 1322
rect -17 1288 17 1322
rect 51 1288 85 1322
rect 119 1288 153 1322
rect 187 1288 221 1322
rect 255 1288 289 1322
rect -415 1173 -381 1207
rect -415 1105 -381 1139
rect -415 1037 -381 1071
rect -415 969 -381 1003
rect -415 901 -381 935
rect -415 833 -381 867
rect -415 765 -381 799
rect -415 697 -381 731
rect -415 629 -381 663
rect -415 561 -381 595
rect -415 493 -381 527
rect -415 425 -381 459
rect -415 357 -381 391
rect -415 289 -381 323
rect -415 221 -381 255
rect -415 153 -381 187
rect -415 85 -381 119
rect -415 17 -381 51
rect -415 -51 -381 -17
rect -415 -119 -381 -85
rect -415 -187 -381 -153
rect -415 -255 -381 -221
rect -415 -323 -381 -289
rect -415 -391 -381 -357
rect -415 -459 -381 -425
rect -415 -527 -381 -493
rect -415 -595 -381 -561
rect -415 -663 -381 -629
rect -415 -731 -381 -697
rect -415 -799 -381 -765
rect -415 -867 -381 -833
rect -415 -935 -381 -901
rect -415 -1003 -381 -969
rect -415 -1071 -381 -1037
rect -415 -1139 -381 -1105
rect -415 -1207 -381 -1173
rect 381 1173 415 1207
rect 381 1105 415 1139
rect 381 1037 415 1071
rect 381 969 415 1003
rect 381 901 415 935
rect 381 833 415 867
rect 381 765 415 799
rect 381 697 415 731
rect 381 629 415 663
rect 381 561 415 595
rect 381 493 415 527
rect 381 425 415 459
rect 381 357 415 391
rect 381 289 415 323
rect 381 221 415 255
rect 381 153 415 187
rect 381 85 415 119
rect 381 17 415 51
rect 381 -51 415 -17
rect 381 -119 415 -85
rect 381 -187 415 -153
rect 381 -255 415 -221
rect 381 -323 415 -289
rect 381 -391 415 -357
rect 381 -459 415 -425
rect 381 -527 415 -493
rect 381 -595 415 -561
rect 381 -663 415 -629
rect 381 -731 415 -697
rect 381 -799 415 -765
rect 381 -867 415 -833
rect 381 -935 415 -901
rect 381 -1003 415 -969
rect 381 -1071 415 -1037
rect 381 -1139 415 -1105
rect 381 -1207 415 -1173
rect -289 -1322 -255 -1288
rect -221 -1322 -187 -1288
rect -153 -1322 -119 -1288
rect -85 -1322 -51 -1288
rect -17 -1322 17 -1288
rect 51 -1322 85 -1288
rect 119 -1322 153 -1288
rect 187 -1322 221 -1288
rect 255 -1322 289 -1288
<< xpolycontact >>
rect -285 760 285 1192
rect -285 -1192 285 -760
<< ppolyres >>
rect -285 -760 285 760
<< locali >>
rect -415 1288 -289 1322
rect -255 1288 -221 1322
rect -187 1288 -153 1322
rect -119 1288 -85 1322
rect -51 1288 -17 1322
rect 17 1288 51 1322
rect 85 1288 119 1322
rect 153 1288 187 1322
rect 221 1288 255 1322
rect 289 1288 415 1322
rect -415 1207 -381 1288
rect 381 1207 415 1288
rect -415 1139 -381 1173
rect -415 1071 -381 1105
rect -415 1003 -381 1037
rect -415 935 -381 969
rect -415 867 -381 901
rect -415 799 -381 833
rect -415 731 -381 765
rect 381 1139 415 1173
rect 381 1071 415 1105
rect 381 1003 415 1037
rect 381 935 415 969
rect 381 867 415 901
rect 381 799 415 833
rect -415 663 -381 697
rect -415 595 -381 629
rect -415 527 -381 561
rect -415 459 -381 493
rect -415 391 -381 425
rect -415 323 -381 357
rect -415 255 -381 289
rect -415 187 -381 221
rect -415 119 -381 153
rect -415 51 -381 85
rect -415 -17 -381 17
rect -415 -85 -381 -51
rect -415 -153 -381 -119
rect -415 -221 -381 -187
rect -415 -289 -381 -255
rect -415 -357 -381 -323
rect -415 -425 -381 -391
rect -415 -493 -381 -459
rect -415 -561 -381 -527
rect -415 -629 -381 -595
rect -415 -697 -381 -663
rect -415 -765 -381 -731
rect 381 731 415 765
rect 381 663 415 697
rect 381 595 415 629
rect 381 527 415 561
rect 381 459 415 493
rect 381 391 415 425
rect 381 323 415 357
rect 381 255 415 289
rect 381 187 415 221
rect 381 119 415 153
rect 381 51 415 85
rect 381 -17 415 17
rect 381 -85 415 -51
rect 381 -153 415 -119
rect 381 -221 415 -187
rect 381 -289 415 -255
rect 381 -357 415 -323
rect 381 -425 415 -391
rect 381 -493 415 -459
rect 381 -561 415 -527
rect 381 -629 415 -595
rect 381 -697 415 -663
rect -415 -833 -381 -799
rect -415 -901 -381 -867
rect -415 -969 -381 -935
rect -415 -1037 -381 -1003
rect -415 -1105 -381 -1071
rect -415 -1173 -381 -1139
rect 381 -765 415 -731
rect 381 -833 415 -799
rect 381 -901 415 -867
rect 381 -969 415 -935
rect 381 -1037 415 -1003
rect 381 -1105 415 -1071
rect 381 -1173 415 -1139
rect -415 -1288 -381 -1207
rect 381 -1288 415 -1207
rect -415 -1322 -289 -1288
rect -255 -1322 -221 -1288
rect -187 -1322 -153 -1288
rect -119 -1322 -85 -1288
rect -51 -1322 -17 -1288
rect 17 -1322 51 -1288
rect 85 -1322 119 -1288
rect 153 -1322 187 -1288
rect 221 -1322 255 -1288
rect 289 -1322 415 -1288
<< viali >>
rect -269 778 269 1172
rect -269 -1173 269 -779
<< metal1 >>
rect -281 1172 281 1180
rect -281 778 -269 1172
rect 269 778 281 1172
rect -281 771 281 778
rect -281 -779 281 -771
rect -281 -1173 -269 -779
rect 269 -1173 281 -779
rect -281 -1180 281 -1173
<< properties >>
string FIXED_BBOX -398 -1305 398 1305
<< end >>
