magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -297 10902 297 10988
rect -297 -10902 -211 10902
rect 211 -10902 297 10902
rect -297 -10988 297 -10902
<< psubdiff >>
rect -271 10928 -153 10962
rect -119 10928 -85 10962
rect -51 10928 -17 10962
rect 17 10928 51 10962
rect 85 10928 119 10962
rect 153 10928 271 10962
rect -271 -10928 -237 10928
rect 237 -10928 271 10928
rect -271 -10962 -153 -10928
rect -119 -10962 -85 -10928
rect -51 -10962 -17 -10928
rect 17 -10962 51 -10928
rect 85 -10962 119 -10928
rect 153 -10962 271 -10928
<< psubdiffcont >>
rect -153 10928 -119 10962
rect -85 10928 -51 10962
rect -17 10928 17 10962
rect 51 10928 85 10962
rect 119 10928 153 10962
rect -153 -10962 -119 -10928
rect -85 -10962 -51 -10928
rect -17 -10962 17 -10928
rect 51 -10962 85 -10928
rect 119 -10962 153 -10928
<< xpolycontact >>
rect -141 10400 141 10832
rect -141 -10832 141 -10400
<< ppolyres >>
rect -141 -10400 141 10400
<< locali >>
rect -271 10928 -153 10962
rect -119 10928 -85 10962
rect -51 10928 -17 10962
rect 17 10928 51 10962
rect 85 10928 119 10962
rect 153 10928 271 10962
rect -271 -10928 -237 10928
rect 237 -10928 271 10928
rect -271 -10962 -153 -10928
rect -119 -10962 -85 -10928
rect -51 -10962 -17 -10928
rect 17 -10962 51 -10928
rect 85 -10962 119 -10928
rect 153 -10962 271 -10928
<< viali >>
rect -125 10418 125 10812
rect -125 -10813 125 -10419
<< metal1 >>
rect -131 10812 131 10826
rect -131 10418 -125 10812
rect 125 10418 131 10812
rect -131 10405 131 10418
rect -131 -10419 131 -10405
rect -131 -10813 -125 -10419
rect 125 -10813 131 -10419
rect -131 -10826 131 -10813
<< properties >>
string FIXED_BBOX -254 -10945 254 10945
<< end >>
