magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -2765 172 -2707 178
rect -2573 172 -2515 178
rect -2381 172 -2323 178
rect -2189 172 -2131 178
rect -1997 172 -1939 178
rect -1805 172 -1747 178
rect -1613 172 -1555 178
rect -1421 172 -1363 178
rect -1229 172 -1171 178
rect -1037 172 -979 178
rect -845 172 -787 178
rect -653 172 -595 178
rect -461 172 -403 178
rect -269 172 -211 178
rect -77 172 -19 178
rect 115 172 173 178
rect 307 172 365 178
rect 499 172 557 178
rect 691 172 749 178
rect 883 172 941 178
rect 1075 172 1133 178
rect 1267 172 1325 178
rect 1459 172 1517 178
rect 1651 172 1709 178
rect 1843 172 1901 178
rect 2035 172 2093 178
rect 2227 172 2285 178
rect 2419 172 2477 178
rect 2611 172 2669 178
rect 2803 172 2861 178
rect -2765 138 -2753 172
rect -2573 138 -2561 172
rect -2381 138 -2369 172
rect -2189 138 -2177 172
rect -1997 138 -1985 172
rect -1805 138 -1793 172
rect -1613 138 -1601 172
rect -1421 138 -1409 172
rect -1229 138 -1217 172
rect -1037 138 -1025 172
rect -845 138 -833 172
rect -653 138 -641 172
rect -461 138 -449 172
rect -269 138 -257 172
rect -77 138 -65 172
rect 115 138 127 172
rect 307 138 319 172
rect 499 138 511 172
rect 691 138 703 172
rect 883 138 895 172
rect 1075 138 1087 172
rect 1267 138 1279 172
rect 1459 138 1471 172
rect 1651 138 1663 172
rect 1843 138 1855 172
rect 2035 138 2047 172
rect 2227 138 2239 172
rect 2419 138 2431 172
rect 2611 138 2623 172
rect 2803 138 2815 172
rect -2765 132 -2707 138
rect -2573 132 -2515 138
rect -2381 132 -2323 138
rect -2189 132 -2131 138
rect -1997 132 -1939 138
rect -1805 132 -1747 138
rect -1613 132 -1555 138
rect -1421 132 -1363 138
rect -1229 132 -1171 138
rect -1037 132 -979 138
rect -845 132 -787 138
rect -653 132 -595 138
rect -461 132 -403 138
rect -269 132 -211 138
rect -77 132 -19 138
rect 115 132 173 138
rect 307 132 365 138
rect 499 132 557 138
rect 691 132 749 138
rect 883 132 941 138
rect 1075 132 1133 138
rect 1267 132 1325 138
rect 1459 132 1517 138
rect 1651 132 1709 138
rect 1843 132 1901 138
rect 2035 132 2093 138
rect 2227 132 2285 138
rect 2419 132 2477 138
rect 2611 132 2669 138
rect 2803 132 2861 138
rect -2861 -138 -2803 -132
rect -2669 -138 -2611 -132
rect -2477 -138 -2419 -132
rect -2285 -138 -2227 -132
rect -2093 -138 -2035 -132
rect -1901 -138 -1843 -132
rect -1709 -138 -1651 -132
rect -1517 -138 -1459 -132
rect -1325 -138 -1267 -132
rect -1133 -138 -1075 -132
rect -941 -138 -883 -132
rect -749 -138 -691 -132
rect -557 -138 -499 -132
rect -365 -138 -307 -132
rect -173 -138 -115 -132
rect 19 -138 77 -132
rect 211 -138 269 -132
rect 403 -138 461 -132
rect 595 -138 653 -132
rect 787 -138 845 -132
rect 979 -138 1037 -132
rect 1171 -138 1229 -132
rect 1363 -138 1421 -132
rect 1555 -138 1613 -132
rect 1747 -138 1805 -132
rect 1939 -138 1997 -132
rect 2131 -138 2189 -132
rect 2323 -138 2381 -132
rect 2515 -138 2573 -132
rect 2707 -138 2765 -132
rect -2861 -172 -2849 -138
rect -2669 -172 -2657 -138
rect -2477 -172 -2465 -138
rect -2285 -172 -2273 -138
rect -2093 -172 -2081 -138
rect -1901 -172 -1889 -138
rect -1709 -172 -1697 -138
rect -1517 -172 -1505 -138
rect -1325 -172 -1313 -138
rect -1133 -172 -1121 -138
rect -941 -172 -929 -138
rect -749 -172 -737 -138
rect -557 -172 -545 -138
rect -365 -172 -353 -138
rect -173 -172 -161 -138
rect 19 -172 31 -138
rect 211 -172 223 -138
rect 403 -172 415 -138
rect 595 -172 607 -138
rect 787 -172 799 -138
rect 979 -172 991 -138
rect 1171 -172 1183 -138
rect 1363 -172 1375 -138
rect 1555 -172 1567 -138
rect 1747 -172 1759 -138
rect 1939 -172 1951 -138
rect 2131 -172 2143 -138
rect 2323 -172 2335 -138
rect 2515 -172 2527 -138
rect 2707 -172 2719 -138
rect -2861 -178 -2803 -172
rect -2669 -178 -2611 -172
rect -2477 -178 -2419 -172
rect -2285 -178 -2227 -172
rect -2093 -178 -2035 -172
rect -1901 -178 -1843 -172
rect -1709 -178 -1651 -172
rect -1517 -178 -1459 -172
rect -1325 -178 -1267 -172
rect -1133 -178 -1075 -172
rect -941 -178 -883 -172
rect -749 -178 -691 -172
rect -557 -178 -499 -172
rect -365 -178 -307 -172
rect -173 -178 -115 -172
rect 19 -178 77 -172
rect 211 -178 269 -172
rect 403 -178 461 -172
rect 595 -178 653 -172
rect 787 -178 845 -172
rect 979 -178 1037 -172
rect 1171 -178 1229 -172
rect 1363 -178 1421 -172
rect 1555 -178 1613 -172
rect 1747 -178 1805 -172
rect 1939 -178 1997 -172
rect 2131 -178 2189 -172
rect 2323 -178 2381 -172
rect 2515 -178 2573 -172
rect 2707 -178 2765 -172
<< pwell >>
rect -3037 -300 3037 300
<< nmoslvt >>
rect -2847 -100 -2817 100
rect -2751 -100 -2721 100
rect -2655 -100 -2625 100
rect -2559 -100 -2529 100
rect -2463 -100 -2433 100
rect -2367 -100 -2337 100
rect -2271 -100 -2241 100
rect -2175 -100 -2145 100
rect -2079 -100 -2049 100
rect -1983 -100 -1953 100
rect -1887 -100 -1857 100
rect -1791 -100 -1761 100
rect -1695 -100 -1665 100
rect -1599 -100 -1569 100
rect -1503 -100 -1473 100
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
rect 1473 -100 1503 100
rect 1569 -100 1599 100
rect 1665 -100 1695 100
rect 1761 -100 1791 100
rect 1857 -100 1887 100
rect 1953 -100 1983 100
rect 2049 -100 2079 100
rect 2145 -100 2175 100
rect 2241 -100 2271 100
rect 2337 -100 2367 100
rect 2433 -100 2463 100
rect 2529 -100 2559 100
rect 2625 -100 2655 100
rect 2721 -100 2751 100
rect 2817 -100 2847 100
<< ndiff >>
rect -2909 85 -2847 100
rect -2909 51 -2897 85
rect -2863 51 -2847 85
rect -2909 17 -2847 51
rect -2909 -17 -2897 17
rect -2863 -17 -2847 17
rect -2909 -51 -2847 -17
rect -2909 -85 -2897 -51
rect -2863 -85 -2847 -51
rect -2909 -100 -2847 -85
rect -2817 85 -2751 100
rect -2817 51 -2801 85
rect -2767 51 -2751 85
rect -2817 17 -2751 51
rect -2817 -17 -2801 17
rect -2767 -17 -2751 17
rect -2817 -51 -2751 -17
rect -2817 -85 -2801 -51
rect -2767 -85 -2751 -51
rect -2817 -100 -2751 -85
rect -2721 85 -2655 100
rect -2721 51 -2705 85
rect -2671 51 -2655 85
rect -2721 17 -2655 51
rect -2721 -17 -2705 17
rect -2671 -17 -2655 17
rect -2721 -51 -2655 -17
rect -2721 -85 -2705 -51
rect -2671 -85 -2655 -51
rect -2721 -100 -2655 -85
rect -2625 85 -2559 100
rect -2625 51 -2609 85
rect -2575 51 -2559 85
rect -2625 17 -2559 51
rect -2625 -17 -2609 17
rect -2575 -17 -2559 17
rect -2625 -51 -2559 -17
rect -2625 -85 -2609 -51
rect -2575 -85 -2559 -51
rect -2625 -100 -2559 -85
rect -2529 85 -2463 100
rect -2529 51 -2513 85
rect -2479 51 -2463 85
rect -2529 17 -2463 51
rect -2529 -17 -2513 17
rect -2479 -17 -2463 17
rect -2529 -51 -2463 -17
rect -2529 -85 -2513 -51
rect -2479 -85 -2463 -51
rect -2529 -100 -2463 -85
rect -2433 85 -2367 100
rect -2433 51 -2417 85
rect -2383 51 -2367 85
rect -2433 17 -2367 51
rect -2433 -17 -2417 17
rect -2383 -17 -2367 17
rect -2433 -51 -2367 -17
rect -2433 -85 -2417 -51
rect -2383 -85 -2367 -51
rect -2433 -100 -2367 -85
rect -2337 85 -2271 100
rect -2337 51 -2321 85
rect -2287 51 -2271 85
rect -2337 17 -2271 51
rect -2337 -17 -2321 17
rect -2287 -17 -2271 17
rect -2337 -51 -2271 -17
rect -2337 -85 -2321 -51
rect -2287 -85 -2271 -51
rect -2337 -100 -2271 -85
rect -2241 85 -2175 100
rect -2241 51 -2225 85
rect -2191 51 -2175 85
rect -2241 17 -2175 51
rect -2241 -17 -2225 17
rect -2191 -17 -2175 17
rect -2241 -51 -2175 -17
rect -2241 -85 -2225 -51
rect -2191 -85 -2175 -51
rect -2241 -100 -2175 -85
rect -2145 85 -2079 100
rect -2145 51 -2129 85
rect -2095 51 -2079 85
rect -2145 17 -2079 51
rect -2145 -17 -2129 17
rect -2095 -17 -2079 17
rect -2145 -51 -2079 -17
rect -2145 -85 -2129 -51
rect -2095 -85 -2079 -51
rect -2145 -100 -2079 -85
rect -2049 85 -1983 100
rect -2049 51 -2033 85
rect -1999 51 -1983 85
rect -2049 17 -1983 51
rect -2049 -17 -2033 17
rect -1999 -17 -1983 17
rect -2049 -51 -1983 -17
rect -2049 -85 -2033 -51
rect -1999 -85 -1983 -51
rect -2049 -100 -1983 -85
rect -1953 85 -1887 100
rect -1953 51 -1937 85
rect -1903 51 -1887 85
rect -1953 17 -1887 51
rect -1953 -17 -1937 17
rect -1903 -17 -1887 17
rect -1953 -51 -1887 -17
rect -1953 -85 -1937 -51
rect -1903 -85 -1887 -51
rect -1953 -100 -1887 -85
rect -1857 85 -1791 100
rect -1857 51 -1841 85
rect -1807 51 -1791 85
rect -1857 17 -1791 51
rect -1857 -17 -1841 17
rect -1807 -17 -1791 17
rect -1857 -51 -1791 -17
rect -1857 -85 -1841 -51
rect -1807 -85 -1791 -51
rect -1857 -100 -1791 -85
rect -1761 85 -1695 100
rect -1761 51 -1745 85
rect -1711 51 -1695 85
rect -1761 17 -1695 51
rect -1761 -17 -1745 17
rect -1711 -17 -1695 17
rect -1761 -51 -1695 -17
rect -1761 -85 -1745 -51
rect -1711 -85 -1695 -51
rect -1761 -100 -1695 -85
rect -1665 85 -1599 100
rect -1665 51 -1649 85
rect -1615 51 -1599 85
rect -1665 17 -1599 51
rect -1665 -17 -1649 17
rect -1615 -17 -1599 17
rect -1665 -51 -1599 -17
rect -1665 -85 -1649 -51
rect -1615 -85 -1599 -51
rect -1665 -100 -1599 -85
rect -1569 85 -1503 100
rect -1569 51 -1553 85
rect -1519 51 -1503 85
rect -1569 17 -1503 51
rect -1569 -17 -1553 17
rect -1519 -17 -1503 17
rect -1569 -51 -1503 -17
rect -1569 -85 -1553 -51
rect -1519 -85 -1503 -51
rect -1569 -100 -1503 -85
rect -1473 85 -1407 100
rect -1473 51 -1457 85
rect -1423 51 -1407 85
rect -1473 17 -1407 51
rect -1473 -17 -1457 17
rect -1423 -17 -1407 17
rect -1473 -51 -1407 -17
rect -1473 -85 -1457 -51
rect -1423 -85 -1407 -51
rect -1473 -100 -1407 -85
rect -1377 85 -1311 100
rect -1377 51 -1361 85
rect -1327 51 -1311 85
rect -1377 17 -1311 51
rect -1377 -17 -1361 17
rect -1327 -17 -1311 17
rect -1377 -51 -1311 -17
rect -1377 -85 -1361 -51
rect -1327 -85 -1311 -51
rect -1377 -100 -1311 -85
rect -1281 85 -1215 100
rect -1281 51 -1265 85
rect -1231 51 -1215 85
rect -1281 17 -1215 51
rect -1281 -17 -1265 17
rect -1231 -17 -1215 17
rect -1281 -51 -1215 -17
rect -1281 -85 -1265 -51
rect -1231 -85 -1215 -51
rect -1281 -100 -1215 -85
rect -1185 85 -1119 100
rect -1185 51 -1169 85
rect -1135 51 -1119 85
rect -1185 17 -1119 51
rect -1185 -17 -1169 17
rect -1135 -17 -1119 17
rect -1185 -51 -1119 -17
rect -1185 -85 -1169 -51
rect -1135 -85 -1119 -51
rect -1185 -100 -1119 -85
rect -1089 85 -1023 100
rect -1089 51 -1073 85
rect -1039 51 -1023 85
rect -1089 17 -1023 51
rect -1089 -17 -1073 17
rect -1039 -17 -1023 17
rect -1089 -51 -1023 -17
rect -1089 -85 -1073 -51
rect -1039 -85 -1023 -51
rect -1089 -100 -1023 -85
rect -993 85 -927 100
rect -993 51 -977 85
rect -943 51 -927 85
rect -993 17 -927 51
rect -993 -17 -977 17
rect -943 -17 -927 17
rect -993 -51 -927 -17
rect -993 -85 -977 -51
rect -943 -85 -927 -51
rect -993 -100 -927 -85
rect -897 85 -831 100
rect -897 51 -881 85
rect -847 51 -831 85
rect -897 17 -831 51
rect -897 -17 -881 17
rect -847 -17 -831 17
rect -897 -51 -831 -17
rect -897 -85 -881 -51
rect -847 -85 -831 -51
rect -897 -100 -831 -85
rect -801 85 -735 100
rect -801 51 -785 85
rect -751 51 -735 85
rect -801 17 -735 51
rect -801 -17 -785 17
rect -751 -17 -735 17
rect -801 -51 -735 -17
rect -801 -85 -785 -51
rect -751 -85 -735 -51
rect -801 -100 -735 -85
rect -705 85 -639 100
rect -705 51 -689 85
rect -655 51 -639 85
rect -705 17 -639 51
rect -705 -17 -689 17
rect -655 -17 -639 17
rect -705 -51 -639 -17
rect -705 -85 -689 -51
rect -655 -85 -639 -51
rect -705 -100 -639 -85
rect -609 85 -543 100
rect -609 51 -593 85
rect -559 51 -543 85
rect -609 17 -543 51
rect -609 -17 -593 17
rect -559 -17 -543 17
rect -609 -51 -543 -17
rect -609 -85 -593 -51
rect -559 -85 -543 -51
rect -609 -100 -543 -85
rect -513 85 -447 100
rect -513 51 -497 85
rect -463 51 -447 85
rect -513 17 -447 51
rect -513 -17 -497 17
rect -463 -17 -447 17
rect -513 -51 -447 -17
rect -513 -85 -497 -51
rect -463 -85 -447 -51
rect -513 -100 -447 -85
rect -417 85 -351 100
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -100 -351 -85
rect -321 85 -255 100
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 321 100
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -100 321 -85
rect 351 85 417 100
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -100 417 -85
rect 447 85 513 100
rect 447 51 463 85
rect 497 51 513 85
rect 447 17 513 51
rect 447 -17 463 17
rect 497 -17 513 17
rect 447 -51 513 -17
rect 447 -85 463 -51
rect 497 -85 513 -51
rect 447 -100 513 -85
rect 543 85 609 100
rect 543 51 559 85
rect 593 51 609 85
rect 543 17 609 51
rect 543 -17 559 17
rect 593 -17 609 17
rect 543 -51 609 -17
rect 543 -85 559 -51
rect 593 -85 609 -51
rect 543 -100 609 -85
rect 639 85 705 100
rect 639 51 655 85
rect 689 51 705 85
rect 639 17 705 51
rect 639 -17 655 17
rect 689 -17 705 17
rect 639 -51 705 -17
rect 639 -85 655 -51
rect 689 -85 705 -51
rect 639 -100 705 -85
rect 735 85 801 100
rect 735 51 751 85
rect 785 51 801 85
rect 735 17 801 51
rect 735 -17 751 17
rect 785 -17 801 17
rect 735 -51 801 -17
rect 735 -85 751 -51
rect 785 -85 801 -51
rect 735 -100 801 -85
rect 831 85 897 100
rect 831 51 847 85
rect 881 51 897 85
rect 831 17 897 51
rect 831 -17 847 17
rect 881 -17 897 17
rect 831 -51 897 -17
rect 831 -85 847 -51
rect 881 -85 897 -51
rect 831 -100 897 -85
rect 927 85 993 100
rect 927 51 943 85
rect 977 51 993 85
rect 927 17 993 51
rect 927 -17 943 17
rect 977 -17 993 17
rect 927 -51 993 -17
rect 927 -85 943 -51
rect 977 -85 993 -51
rect 927 -100 993 -85
rect 1023 85 1089 100
rect 1023 51 1039 85
rect 1073 51 1089 85
rect 1023 17 1089 51
rect 1023 -17 1039 17
rect 1073 -17 1089 17
rect 1023 -51 1089 -17
rect 1023 -85 1039 -51
rect 1073 -85 1089 -51
rect 1023 -100 1089 -85
rect 1119 85 1185 100
rect 1119 51 1135 85
rect 1169 51 1185 85
rect 1119 17 1185 51
rect 1119 -17 1135 17
rect 1169 -17 1185 17
rect 1119 -51 1185 -17
rect 1119 -85 1135 -51
rect 1169 -85 1185 -51
rect 1119 -100 1185 -85
rect 1215 85 1281 100
rect 1215 51 1231 85
rect 1265 51 1281 85
rect 1215 17 1281 51
rect 1215 -17 1231 17
rect 1265 -17 1281 17
rect 1215 -51 1281 -17
rect 1215 -85 1231 -51
rect 1265 -85 1281 -51
rect 1215 -100 1281 -85
rect 1311 85 1377 100
rect 1311 51 1327 85
rect 1361 51 1377 85
rect 1311 17 1377 51
rect 1311 -17 1327 17
rect 1361 -17 1377 17
rect 1311 -51 1377 -17
rect 1311 -85 1327 -51
rect 1361 -85 1377 -51
rect 1311 -100 1377 -85
rect 1407 85 1473 100
rect 1407 51 1423 85
rect 1457 51 1473 85
rect 1407 17 1473 51
rect 1407 -17 1423 17
rect 1457 -17 1473 17
rect 1407 -51 1473 -17
rect 1407 -85 1423 -51
rect 1457 -85 1473 -51
rect 1407 -100 1473 -85
rect 1503 85 1569 100
rect 1503 51 1519 85
rect 1553 51 1569 85
rect 1503 17 1569 51
rect 1503 -17 1519 17
rect 1553 -17 1569 17
rect 1503 -51 1569 -17
rect 1503 -85 1519 -51
rect 1553 -85 1569 -51
rect 1503 -100 1569 -85
rect 1599 85 1665 100
rect 1599 51 1615 85
rect 1649 51 1665 85
rect 1599 17 1665 51
rect 1599 -17 1615 17
rect 1649 -17 1665 17
rect 1599 -51 1665 -17
rect 1599 -85 1615 -51
rect 1649 -85 1665 -51
rect 1599 -100 1665 -85
rect 1695 85 1761 100
rect 1695 51 1711 85
rect 1745 51 1761 85
rect 1695 17 1761 51
rect 1695 -17 1711 17
rect 1745 -17 1761 17
rect 1695 -51 1761 -17
rect 1695 -85 1711 -51
rect 1745 -85 1761 -51
rect 1695 -100 1761 -85
rect 1791 85 1857 100
rect 1791 51 1807 85
rect 1841 51 1857 85
rect 1791 17 1857 51
rect 1791 -17 1807 17
rect 1841 -17 1857 17
rect 1791 -51 1857 -17
rect 1791 -85 1807 -51
rect 1841 -85 1857 -51
rect 1791 -100 1857 -85
rect 1887 85 1953 100
rect 1887 51 1903 85
rect 1937 51 1953 85
rect 1887 17 1953 51
rect 1887 -17 1903 17
rect 1937 -17 1953 17
rect 1887 -51 1953 -17
rect 1887 -85 1903 -51
rect 1937 -85 1953 -51
rect 1887 -100 1953 -85
rect 1983 85 2049 100
rect 1983 51 1999 85
rect 2033 51 2049 85
rect 1983 17 2049 51
rect 1983 -17 1999 17
rect 2033 -17 2049 17
rect 1983 -51 2049 -17
rect 1983 -85 1999 -51
rect 2033 -85 2049 -51
rect 1983 -100 2049 -85
rect 2079 85 2145 100
rect 2079 51 2095 85
rect 2129 51 2145 85
rect 2079 17 2145 51
rect 2079 -17 2095 17
rect 2129 -17 2145 17
rect 2079 -51 2145 -17
rect 2079 -85 2095 -51
rect 2129 -85 2145 -51
rect 2079 -100 2145 -85
rect 2175 85 2241 100
rect 2175 51 2191 85
rect 2225 51 2241 85
rect 2175 17 2241 51
rect 2175 -17 2191 17
rect 2225 -17 2241 17
rect 2175 -51 2241 -17
rect 2175 -85 2191 -51
rect 2225 -85 2241 -51
rect 2175 -100 2241 -85
rect 2271 85 2337 100
rect 2271 51 2287 85
rect 2321 51 2337 85
rect 2271 17 2337 51
rect 2271 -17 2287 17
rect 2321 -17 2337 17
rect 2271 -51 2337 -17
rect 2271 -85 2287 -51
rect 2321 -85 2337 -51
rect 2271 -100 2337 -85
rect 2367 85 2433 100
rect 2367 51 2383 85
rect 2417 51 2433 85
rect 2367 17 2433 51
rect 2367 -17 2383 17
rect 2417 -17 2433 17
rect 2367 -51 2433 -17
rect 2367 -85 2383 -51
rect 2417 -85 2433 -51
rect 2367 -100 2433 -85
rect 2463 85 2529 100
rect 2463 51 2479 85
rect 2513 51 2529 85
rect 2463 17 2529 51
rect 2463 -17 2479 17
rect 2513 -17 2529 17
rect 2463 -51 2529 -17
rect 2463 -85 2479 -51
rect 2513 -85 2529 -51
rect 2463 -100 2529 -85
rect 2559 85 2625 100
rect 2559 51 2575 85
rect 2609 51 2625 85
rect 2559 17 2625 51
rect 2559 -17 2575 17
rect 2609 -17 2625 17
rect 2559 -51 2625 -17
rect 2559 -85 2575 -51
rect 2609 -85 2625 -51
rect 2559 -100 2625 -85
rect 2655 85 2721 100
rect 2655 51 2671 85
rect 2705 51 2721 85
rect 2655 17 2721 51
rect 2655 -17 2671 17
rect 2705 -17 2721 17
rect 2655 -51 2721 -17
rect 2655 -85 2671 -51
rect 2705 -85 2721 -51
rect 2655 -100 2721 -85
rect 2751 85 2817 100
rect 2751 51 2767 85
rect 2801 51 2817 85
rect 2751 17 2817 51
rect 2751 -17 2767 17
rect 2801 -17 2817 17
rect 2751 -51 2817 -17
rect 2751 -85 2767 -51
rect 2801 -85 2817 -51
rect 2751 -100 2817 -85
rect 2847 85 2909 100
rect 2847 51 2863 85
rect 2897 51 2909 85
rect 2847 17 2909 51
rect 2847 -17 2863 17
rect 2897 -17 2909 17
rect 2847 -51 2909 -17
rect 2847 -85 2863 -51
rect 2897 -85 2909 -51
rect 2847 -100 2909 -85
<< ndiffc >>
rect -2897 51 -2863 85
rect -2897 -17 -2863 17
rect -2897 -85 -2863 -51
rect -2801 51 -2767 85
rect -2801 -17 -2767 17
rect -2801 -85 -2767 -51
rect -2705 51 -2671 85
rect -2705 -17 -2671 17
rect -2705 -85 -2671 -51
rect -2609 51 -2575 85
rect -2609 -17 -2575 17
rect -2609 -85 -2575 -51
rect -2513 51 -2479 85
rect -2513 -17 -2479 17
rect -2513 -85 -2479 -51
rect -2417 51 -2383 85
rect -2417 -17 -2383 17
rect -2417 -85 -2383 -51
rect -2321 51 -2287 85
rect -2321 -17 -2287 17
rect -2321 -85 -2287 -51
rect -2225 51 -2191 85
rect -2225 -17 -2191 17
rect -2225 -85 -2191 -51
rect -2129 51 -2095 85
rect -2129 -17 -2095 17
rect -2129 -85 -2095 -51
rect -2033 51 -1999 85
rect -2033 -17 -1999 17
rect -2033 -85 -1999 -51
rect -1937 51 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -51
rect -1841 51 -1807 85
rect -1841 -17 -1807 17
rect -1841 -85 -1807 -51
rect -1745 51 -1711 85
rect -1745 -17 -1711 17
rect -1745 -85 -1711 -51
rect -1649 51 -1615 85
rect -1649 -17 -1615 17
rect -1649 -85 -1615 -51
rect -1553 51 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -51
rect -1457 51 -1423 85
rect -1457 -17 -1423 17
rect -1457 -85 -1423 -51
rect -1361 51 -1327 85
rect -1361 -17 -1327 17
rect -1361 -85 -1327 -51
rect -1265 51 -1231 85
rect -1265 -17 -1231 17
rect -1265 -85 -1231 -51
rect -1169 51 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -51
rect -1073 51 -1039 85
rect -1073 -17 -1039 17
rect -1073 -85 -1039 -51
rect -977 51 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -51
rect -881 51 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -51
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -689 51 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -51
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 655 51 689 85
rect 655 -17 689 17
rect 655 -85 689 -51
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 847 51 881 85
rect 847 -17 881 17
rect 847 -85 881 -51
rect 943 51 977 85
rect 943 -17 977 17
rect 943 -85 977 -51
rect 1039 51 1073 85
rect 1039 -17 1073 17
rect 1039 -85 1073 -51
rect 1135 51 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -51
rect 1231 51 1265 85
rect 1231 -17 1265 17
rect 1231 -85 1265 -51
rect 1327 51 1361 85
rect 1327 -17 1361 17
rect 1327 -85 1361 -51
rect 1423 51 1457 85
rect 1423 -17 1457 17
rect 1423 -85 1457 -51
rect 1519 51 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -51
rect 1615 51 1649 85
rect 1615 -17 1649 17
rect 1615 -85 1649 -51
rect 1711 51 1745 85
rect 1711 -17 1745 17
rect 1711 -85 1745 -51
rect 1807 51 1841 85
rect 1807 -17 1841 17
rect 1807 -85 1841 -51
rect 1903 51 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -51
rect 1999 51 2033 85
rect 1999 -17 2033 17
rect 1999 -85 2033 -51
rect 2095 51 2129 85
rect 2095 -17 2129 17
rect 2095 -85 2129 -51
rect 2191 51 2225 85
rect 2191 -17 2225 17
rect 2191 -85 2225 -51
rect 2287 51 2321 85
rect 2287 -17 2321 17
rect 2287 -85 2321 -51
rect 2383 51 2417 85
rect 2383 -17 2417 17
rect 2383 -85 2417 -51
rect 2479 51 2513 85
rect 2479 -17 2513 17
rect 2479 -85 2513 -51
rect 2575 51 2609 85
rect 2575 -17 2609 17
rect 2575 -85 2609 -51
rect 2671 51 2705 85
rect 2671 -17 2705 17
rect 2671 -85 2705 -51
rect 2767 51 2801 85
rect 2767 -17 2801 17
rect 2767 -85 2801 -51
rect 2863 51 2897 85
rect 2863 -17 2897 17
rect 2863 -85 2897 -51
<< psubdiff >>
rect -3011 240 -2907 274
rect -2873 240 -2839 274
rect -2805 240 -2771 274
rect -2737 240 -2703 274
rect -2669 240 -2635 274
rect -2601 240 -2567 274
rect -2533 240 -2499 274
rect -2465 240 -2431 274
rect -2397 240 -2363 274
rect -2329 240 -2295 274
rect -2261 240 -2227 274
rect -2193 240 -2159 274
rect -2125 240 -2091 274
rect -2057 240 -2023 274
rect -1989 240 -1955 274
rect -1921 240 -1887 274
rect -1853 240 -1819 274
rect -1785 240 -1751 274
rect -1717 240 -1683 274
rect -1649 240 -1615 274
rect -1581 240 -1547 274
rect -1513 240 -1479 274
rect -1445 240 -1411 274
rect -1377 240 -1343 274
rect -1309 240 -1275 274
rect -1241 240 -1207 274
rect -1173 240 -1139 274
rect -1105 240 -1071 274
rect -1037 240 -1003 274
rect -969 240 -935 274
rect -901 240 -867 274
rect -833 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 833 274
rect 867 240 901 274
rect 935 240 969 274
rect 1003 240 1037 274
rect 1071 240 1105 274
rect 1139 240 1173 274
rect 1207 240 1241 274
rect 1275 240 1309 274
rect 1343 240 1377 274
rect 1411 240 1445 274
rect 1479 240 1513 274
rect 1547 240 1581 274
rect 1615 240 1649 274
rect 1683 240 1717 274
rect 1751 240 1785 274
rect 1819 240 1853 274
rect 1887 240 1921 274
rect 1955 240 1989 274
rect 2023 240 2057 274
rect 2091 240 2125 274
rect 2159 240 2193 274
rect 2227 240 2261 274
rect 2295 240 2329 274
rect 2363 240 2397 274
rect 2431 240 2465 274
rect 2499 240 2533 274
rect 2567 240 2601 274
rect 2635 240 2669 274
rect 2703 240 2737 274
rect 2771 240 2805 274
rect 2839 240 2873 274
rect 2907 240 3011 274
rect -3011 153 -2977 240
rect -3011 85 -2977 119
rect 2977 153 3011 240
rect -3011 17 -2977 51
rect -3011 -51 -2977 -17
rect -3011 -119 -2977 -85
rect 2977 85 3011 119
rect 2977 17 3011 51
rect 2977 -51 3011 -17
rect -3011 -240 -2977 -153
rect 2977 -119 3011 -85
rect 2977 -240 3011 -153
rect -3011 -274 -2907 -240
rect -2873 -274 -2839 -240
rect -2805 -274 -2771 -240
rect -2737 -274 -2703 -240
rect -2669 -274 -2635 -240
rect -2601 -274 -2567 -240
rect -2533 -274 -2499 -240
rect -2465 -274 -2431 -240
rect -2397 -274 -2363 -240
rect -2329 -274 -2295 -240
rect -2261 -274 -2227 -240
rect -2193 -274 -2159 -240
rect -2125 -274 -2091 -240
rect -2057 -274 -2023 -240
rect -1989 -274 -1955 -240
rect -1921 -274 -1887 -240
rect -1853 -274 -1819 -240
rect -1785 -274 -1751 -240
rect -1717 -274 -1683 -240
rect -1649 -274 -1615 -240
rect -1581 -274 -1547 -240
rect -1513 -274 -1479 -240
rect -1445 -274 -1411 -240
rect -1377 -274 -1343 -240
rect -1309 -274 -1275 -240
rect -1241 -274 -1207 -240
rect -1173 -274 -1139 -240
rect -1105 -274 -1071 -240
rect -1037 -274 -1003 -240
rect -969 -274 -935 -240
rect -901 -274 -867 -240
rect -833 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 833 -240
rect 867 -274 901 -240
rect 935 -274 969 -240
rect 1003 -274 1037 -240
rect 1071 -274 1105 -240
rect 1139 -274 1173 -240
rect 1207 -274 1241 -240
rect 1275 -274 1309 -240
rect 1343 -274 1377 -240
rect 1411 -274 1445 -240
rect 1479 -274 1513 -240
rect 1547 -274 1581 -240
rect 1615 -274 1649 -240
rect 1683 -274 1717 -240
rect 1751 -274 1785 -240
rect 1819 -274 1853 -240
rect 1887 -274 1921 -240
rect 1955 -274 1989 -240
rect 2023 -274 2057 -240
rect 2091 -274 2125 -240
rect 2159 -274 2193 -240
rect 2227 -274 2261 -240
rect 2295 -274 2329 -240
rect 2363 -274 2397 -240
rect 2431 -274 2465 -240
rect 2499 -274 2533 -240
rect 2567 -274 2601 -240
rect 2635 -274 2669 -240
rect 2703 -274 2737 -240
rect 2771 -274 2805 -240
rect 2839 -274 2873 -240
rect 2907 -274 3011 -240
<< psubdiffcont >>
rect -2907 240 -2873 274
rect -2839 240 -2805 274
rect -2771 240 -2737 274
rect -2703 240 -2669 274
rect -2635 240 -2601 274
rect -2567 240 -2533 274
rect -2499 240 -2465 274
rect -2431 240 -2397 274
rect -2363 240 -2329 274
rect -2295 240 -2261 274
rect -2227 240 -2193 274
rect -2159 240 -2125 274
rect -2091 240 -2057 274
rect -2023 240 -1989 274
rect -1955 240 -1921 274
rect -1887 240 -1853 274
rect -1819 240 -1785 274
rect -1751 240 -1717 274
rect -1683 240 -1649 274
rect -1615 240 -1581 274
rect -1547 240 -1513 274
rect -1479 240 -1445 274
rect -1411 240 -1377 274
rect -1343 240 -1309 274
rect -1275 240 -1241 274
rect -1207 240 -1173 274
rect -1139 240 -1105 274
rect -1071 240 -1037 274
rect -1003 240 -969 274
rect -935 240 -901 274
rect -867 240 -833 274
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect 833 240 867 274
rect 901 240 935 274
rect 969 240 1003 274
rect 1037 240 1071 274
rect 1105 240 1139 274
rect 1173 240 1207 274
rect 1241 240 1275 274
rect 1309 240 1343 274
rect 1377 240 1411 274
rect 1445 240 1479 274
rect 1513 240 1547 274
rect 1581 240 1615 274
rect 1649 240 1683 274
rect 1717 240 1751 274
rect 1785 240 1819 274
rect 1853 240 1887 274
rect 1921 240 1955 274
rect 1989 240 2023 274
rect 2057 240 2091 274
rect 2125 240 2159 274
rect 2193 240 2227 274
rect 2261 240 2295 274
rect 2329 240 2363 274
rect 2397 240 2431 274
rect 2465 240 2499 274
rect 2533 240 2567 274
rect 2601 240 2635 274
rect 2669 240 2703 274
rect 2737 240 2771 274
rect 2805 240 2839 274
rect 2873 240 2907 274
rect -3011 119 -2977 153
rect 2977 119 3011 153
rect -3011 51 -2977 85
rect -3011 -17 -2977 17
rect -3011 -85 -2977 -51
rect 2977 51 3011 85
rect 2977 -17 3011 17
rect 2977 -85 3011 -51
rect -3011 -153 -2977 -119
rect 2977 -153 3011 -119
rect -2907 -274 -2873 -240
rect -2839 -274 -2805 -240
rect -2771 -274 -2737 -240
rect -2703 -274 -2669 -240
rect -2635 -274 -2601 -240
rect -2567 -274 -2533 -240
rect -2499 -274 -2465 -240
rect -2431 -274 -2397 -240
rect -2363 -274 -2329 -240
rect -2295 -274 -2261 -240
rect -2227 -274 -2193 -240
rect -2159 -274 -2125 -240
rect -2091 -274 -2057 -240
rect -2023 -274 -1989 -240
rect -1955 -274 -1921 -240
rect -1887 -274 -1853 -240
rect -1819 -274 -1785 -240
rect -1751 -274 -1717 -240
rect -1683 -274 -1649 -240
rect -1615 -274 -1581 -240
rect -1547 -274 -1513 -240
rect -1479 -274 -1445 -240
rect -1411 -274 -1377 -240
rect -1343 -274 -1309 -240
rect -1275 -274 -1241 -240
rect -1207 -274 -1173 -240
rect -1139 -274 -1105 -240
rect -1071 -274 -1037 -240
rect -1003 -274 -969 -240
rect -935 -274 -901 -240
rect -867 -274 -833 -240
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
rect 833 -274 867 -240
rect 901 -274 935 -240
rect 969 -274 1003 -240
rect 1037 -274 1071 -240
rect 1105 -274 1139 -240
rect 1173 -274 1207 -240
rect 1241 -274 1275 -240
rect 1309 -274 1343 -240
rect 1377 -274 1411 -240
rect 1445 -274 1479 -240
rect 1513 -274 1547 -240
rect 1581 -274 1615 -240
rect 1649 -274 1683 -240
rect 1717 -274 1751 -240
rect 1785 -274 1819 -240
rect 1853 -274 1887 -240
rect 1921 -274 1955 -240
rect 1989 -274 2023 -240
rect 2057 -274 2091 -240
rect 2125 -274 2159 -240
rect 2193 -274 2227 -240
rect 2261 -274 2295 -240
rect 2329 -274 2363 -240
rect 2397 -274 2431 -240
rect 2465 -274 2499 -240
rect 2533 -274 2567 -240
rect 2601 -274 2635 -240
rect 2669 -274 2703 -240
rect 2737 -274 2771 -240
rect 2805 -274 2839 -240
rect 2873 -274 2907 -240
<< poly >>
rect -2769 172 -2703 188
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2847 100 -2817 126
rect -2769 122 -2703 138
rect -2577 172 -2511 188
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2751 100 -2721 122
rect -2655 100 -2625 126
rect -2577 122 -2511 138
rect -2385 172 -2319 188
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2559 100 -2529 122
rect -2463 100 -2433 126
rect -2385 122 -2319 138
rect -2193 172 -2127 188
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2367 100 -2337 122
rect -2271 100 -2241 126
rect -2193 122 -2127 138
rect -2001 172 -1935 188
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -2175 100 -2145 122
rect -2079 100 -2049 126
rect -2001 122 -1935 138
rect -1809 172 -1743 188
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1983 100 -1953 122
rect -1887 100 -1857 126
rect -1809 122 -1743 138
rect -1617 172 -1551 188
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1791 100 -1761 122
rect -1695 100 -1665 126
rect -1617 122 -1551 138
rect -1425 172 -1359 188
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1599 100 -1569 122
rect -1503 100 -1473 126
rect -1425 122 -1359 138
rect -1233 172 -1167 188
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1407 100 -1377 122
rect -1311 100 -1281 126
rect -1233 122 -1167 138
rect -1041 172 -975 188
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -1215 100 -1185 122
rect -1119 100 -1089 126
rect -1041 122 -975 138
rect -849 172 -783 188
rect -849 138 -833 172
rect -799 138 -783 172
rect -1023 100 -993 122
rect -927 100 -897 126
rect -849 122 -783 138
rect -657 172 -591 188
rect -657 138 -641 172
rect -607 138 -591 172
rect -831 100 -801 122
rect -735 100 -705 126
rect -657 122 -591 138
rect -465 172 -399 188
rect -465 138 -449 172
rect -415 138 -399 172
rect -639 100 -609 122
rect -543 100 -513 126
rect -465 122 -399 138
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -447 100 -417 122
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 495 172 561 188
rect 495 138 511 172
rect 545 138 561 172
rect 321 100 351 122
rect 417 100 447 126
rect 495 122 561 138
rect 687 172 753 188
rect 687 138 703 172
rect 737 138 753 172
rect 513 100 543 122
rect 609 100 639 126
rect 687 122 753 138
rect 879 172 945 188
rect 879 138 895 172
rect 929 138 945 172
rect 705 100 735 122
rect 801 100 831 126
rect 879 122 945 138
rect 1071 172 1137 188
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 897 100 927 122
rect 993 100 1023 126
rect 1071 122 1137 138
rect 1263 172 1329 188
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1089 100 1119 122
rect 1185 100 1215 126
rect 1263 122 1329 138
rect 1455 172 1521 188
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1281 100 1311 122
rect 1377 100 1407 126
rect 1455 122 1521 138
rect 1647 172 1713 188
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1473 100 1503 122
rect 1569 100 1599 126
rect 1647 122 1713 138
rect 1839 172 1905 188
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 1665 100 1695 122
rect 1761 100 1791 126
rect 1839 122 1905 138
rect 2031 172 2097 188
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 1857 100 1887 122
rect 1953 100 1983 126
rect 2031 122 2097 138
rect 2223 172 2289 188
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2049 100 2079 122
rect 2145 100 2175 126
rect 2223 122 2289 138
rect 2415 172 2481 188
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2241 100 2271 122
rect 2337 100 2367 126
rect 2415 122 2481 138
rect 2607 172 2673 188
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2433 100 2463 122
rect 2529 100 2559 126
rect 2607 122 2673 138
rect 2799 172 2865 188
rect 2799 138 2815 172
rect 2849 138 2865 172
rect 2625 100 2655 122
rect 2721 100 2751 126
rect 2799 122 2865 138
rect 2817 100 2847 122
rect -2847 -122 -2817 -100
rect -2865 -138 -2799 -122
rect -2751 -126 -2721 -100
rect -2655 -122 -2625 -100
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2865 -188 -2799 -172
rect -2673 -138 -2607 -122
rect -2559 -126 -2529 -100
rect -2463 -122 -2433 -100
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2673 -188 -2607 -172
rect -2481 -138 -2415 -122
rect -2367 -126 -2337 -100
rect -2271 -122 -2241 -100
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2481 -188 -2415 -172
rect -2289 -138 -2223 -122
rect -2175 -126 -2145 -100
rect -2079 -122 -2049 -100
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2289 -188 -2223 -172
rect -2097 -138 -2031 -122
rect -1983 -126 -1953 -100
rect -1887 -122 -1857 -100
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -2097 -188 -2031 -172
rect -1905 -138 -1839 -122
rect -1791 -126 -1761 -100
rect -1695 -122 -1665 -100
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1905 -188 -1839 -172
rect -1713 -138 -1647 -122
rect -1599 -126 -1569 -100
rect -1503 -122 -1473 -100
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1713 -188 -1647 -172
rect -1521 -138 -1455 -122
rect -1407 -126 -1377 -100
rect -1311 -122 -1281 -100
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1521 -188 -1455 -172
rect -1329 -138 -1263 -122
rect -1215 -126 -1185 -100
rect -1119 -122 -1089 -100
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1329 -188 -1263 -172
rect -1137 -138 -1071 -122
rect -1023 -126 -993 -100
rect -927 -122 -897 -100
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -1137 -188 -1071 -172
rect -945 -138 -879 -122
rect -831 -126 -801 -100
rect -735 -122 -705 -100
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -945 -188 -879 -172
rect -753 -138 -687 -122
rect -639 -126 -609 -100
rect -543 -122 -513 -100
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -753 -188 -687 -172
rect -561 -138 -495 -122
rect -447 -126 -417 -100
rect -351 -122 -321 -100
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -561 -188 -495 -172
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 417 -122 447 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
rect 399 -138 465 -122
rect 513 -126 543 -100
rect 609 -122 639 -100
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 399 -188 465 -172
rect 591 -138 657 -122
rect 705 -126 735 -100
rect 801 -122 831 -100
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 591 -188 657 -172
rect 783 -138 849 -122
rect 897 -126 927 -100
rect 993 -122 1023 -100
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 783 -188 849 -172
rect 975 -138 1041 -122
rect 1089 -126 1119 -100
rect 1185 -122 1215 -100
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 975 -188 1041 -172
rect 1167 -138 1233 -122
rect 1281 -126 1311 -100
rect 1377 -122 1407 -100
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1167 -188 1233 -172
rect 1359 -138 1425 -122
rect 1473 -126 1503 -100
rect 1569 -122 1599 -100
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1359 -188 1425 -172
rect 1551 -138 1617 -122
rect 1665 -126 1695 -100
rect 1761 -122 1791 -100
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1551 -188 1617 -172
rect 1743 -138 1809 -122
rect 1857 -126 1887 -100
rect 1953 -122 1983 -100
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1743 -188 1809 -172
rect 1935 -138 2001 -122
rect 2049 -126 2079 -100
rect 2145 -122 2175 -100
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 1935 -188 2001 -172
rect 2127 -138 2193 -122
rect 2241 -126 2271 -100
rect 2337 -122 2367 -100
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2127 -188 2193 -172
rect 2319 -138 2385 -122
rect 2433 -126 2463 -100
rect 2529 -122 2559 -100
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2319 -188 2385 -172
rect 2511 -138 2577 -122
rect 2625 -126 2655 -100
rect 2721 -122 2751 -100
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2511 -188 2577 -172
rect 2703 -138 2769 -122
rect 2817 -126 2847 -100
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect 2703 -188 2769 -172
<< polycont >>
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
<< locali >>
rect -3011 240 -2907 274
rect -2873 240 -2839 274
rect -2805 240 -2771 274
rect -2737 240 -2703 274
rect -2669 240 -2635 274
rect -2601 240 -2567 274
rect -2533 240 -2499 274
rect -2465 240 -2431 274
rect -2397 240 -2363 274
rect -2329 240 -2295 274
rect -2261 240 -2227 274
rect -2193 240 -2159 274
rect -2125 240 -2091 274
rect -2057 240 -2023 274
rect -1989 240 -1955 274
rect -1921 240 -1887 274
rect -1853 240 -1819 274
rect -1785 240 -1751 274
rect -1717 240 -1683 274
rect -1649 240 -1615 274
rect -1581 240 -1547 274
rect -1513 240 -1479 274
rect -1445 240 -1411 274
rect -1377 240 -1343 274
rect -1309 240 -1275 274
rect -1241 240 -1207 274
rect -1173 240 -1139 274
rect -1105 240 -1071 274
rect -1037 240 -1003 274
rect -969 240 -935 274
rect -901 240 -867 274
rect -833 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 833 274
rect 867 240 901 274
rect 935 240 969 274
rect 1003 240 1037 274
rect 1071 240 1105 274
rect 1139 240 1173 274
rect 1207 240 1241 274
rect 1275 240 1309 274
rect 1343 240 1377 274
rect 1411 240 1445 274
rect 1479 240 1513 274
rect 1547 240 1581 274
rect 1615 240 1649 274
rect 1683 240 1717 274
rect 1751 240 1785 274
rect 1819 240 1853 274
rect 1887 240 1921 274
rect 1955 240 1989 274
rect 2023 240 2057 274
rect 2091 240 2125 274
rect 2159 240 2193 274
rect 2227 240 2261 274
rect 2295 240 2329 274
rect 2363 240 2397 274
rect 2431 240 2465 274
rect 2499 240 2533 274
rect 2567 240 2601 274
rect 2635 240 2669 274
rect 2703 240 2737 274
rect 2771 240 2805 274
rect 2839 240 2873 274
rect 2907 240 3011 274
rect -3011 153 -2977 240
rect -2769 138 -2753 172
rect -2719 138 -2703 172
rect -2577 138 -2561 172
rect -2527 138 -2511 172
rect -2385 138 -2369 172
rect -2335 138 -2319 172
rect -2193 138 -2177 172
rect -2143 138 -2127 172
rect -2001 138 -1985 172
rect -1951 138 -1935 172
rect -1809 138 -1793 172
rect -1759 138 -1743 172
rect -1617 138 -1601 172
rect -1567 138 -1551 172
rect -1425 138 -1409 172
rect -1375 138 -1359 172
rect -1233 138 -1217 172
rect -1183 138 -1167 172
rect -1041 138 -1025 172
rect -991 138 -975 172
rect -849 138 -833 172
rect -799 138 -783 172
rect -657 138 -641 172
rect -607 138 -591 172
rect -465 138 -449 172
rect -415 138 -399 172
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect 495 138 511 172
rect 545 138 561 172
rect 687 138 703 172
rect 737 138 753 172
rect 879 138 895 172
rect 929 138 945 172
rect 1071 138 1087 172
rect 1121 138 1137 172
rect 1263 138 1279 172
rect 1313 138 1329 172
rect 1455 138 1471 172
rect 1505 138 1521 172
rect 1647 138 1663 172
rect 1697 138 1713 172
rect 1839 138 1855 172
rect 1889 138 1905 172
rect 2031 138 2047 172
rect 2081 138 2097 172
rect 2223 138 2239 172
rect 2273 138 2289 172
rect 2415 138 2431 172
rect 2465 138 2481 172
rect 2607 138 2623 172
rect 2657 138 2673 172
rect 2799 138 2815 172
rect 2849 138 2865 172
rect 2977 153 3011 240
rect -3011 85 -2977 119
rect -3011 17 -2977 51
rect -3011 -51 -2977 -17
rect -3011 -119 -2977 -85
rect -2897 85 -2863 104
rect -2897 17 -2863 19
rect -2897 -19 -2863 -17
rect -2897 -104 -2863 -85
rect -2801 85 -2767 104
rect -2801 17 -2767 19
rect -2801 -19 -2767 -17
rect -2801 -104 -2767 -85
rect -2705 85 -2671 104
rect -2705 17 -2671 19
rect -2705 -19 -2671 -17
rect -2705 -104 -2671 -85
rect -2609 85 -2575 104
rect -2609 17 -2575 19
rect -2609 -19 -2575 -17
rect -2609 -104 -2575 -85
rect -2513 85 -2479 104
rect -2513 17 -2479 19
rect -2513 -19 -2479 -17
rect -2513 -104 -2479 -85
rect -2417 85 -2383 104
rect -2417 17 -2383 19
rect -2417 -19 -2383 -17
rect -2417 -104 -2383 -85
rect -2321 85 -2287 104
rect -2321 17 -2287 19
rect -2321 -19 -2287 -17
rect -2321 -104 -2287 -85
rect -2225 85 -2191 104
rect -2225 17 -2191 19
rect -2225 -19 -2191 -17
rect -2225 -104 -2191 -85
rect -2129 85 -2095 104
rect -2129 17 -2095 19
rect -2129 -19 -2095 -17
rect -2129 -104 -2095 -85
rect -2033 85 -1999 104
rect -2033 17 -1999 19
rect -2033 -19 -1999 -17
rect -2033 -104 -1999 -85
rect -1937 85 -1903 104
rect -1937 17 -1903 19
rect -1937 -19 -1903 -17
rect -1937 -104 -1903 -85
rect -1841 85 -1807 104
rect -1841 17 -1807 19
rect -1841 -19 -1807 -17
rect -1841 -104 -1807 -85
rect -1745 85 -1711 104
rect -1745 17 -1711 19
rect -1745 -19 -1711 -17
rect -1745 -104 -1711 -85
rect -1649 85 -1615 104
rect -1649 17 -1615 19
rect -1649 -19 -1615 -17
rect -1649 -104 -1615 -85
rect -1553 85 -1519 104
rect -1553 17 -1519 19
rect -1553 -19 -1519 -17
rect -1553 -104 -1519 -85
rect -1457 85 -1423 104
rect -1457 17 -1423 19
rect -1457 -19 -1423 -17
rect -1457 -104 -1423 -85
rect -1361 85 -1327 104
rect -1361 17 -1327 19
rect -1361 -19 -1327 -17
rect -1361 -104 -1327 -85
rect -1265 85 -1231 104
rect -1265 17 -1231 19
rect -1265 -19 -1231 -17
rect -1265 -104 -1231 -85
rect -1169 85 -1135 104
rect -1169 17 -1135 19
rect -1169 -19 -1135 -17
rect -1169 -104 -1135 -85
rect -1073 85 -1039 104
rect -1073 17 -1039 19
rect -1073 -19 -1039 -17
rect -1073 -104 -1039 -85
rect -977 85 -943 104
rect -977 17 -943 19
rect -977 -19 -943 -17
rect -977 -104 -943 -85
rect -881 85 -847 104
rect -881 17 -847 19
rect -881 -19 -847 -17
rect -881 -104 -847 -85
rect -785 85 -751 104
rect -785 17 -751 19
rect -785 -19 -751 -17
rect -785 -104 -751 -85
rect -689 85 -655 104
rect -689 17 -655 19
rect -689 -19 -655 -17
rect -689 -104 -655 -85
rect -593 85 -559 104
rect -593 17 -559 19
rect -593 -19 -559 -17
rect -593 -104 -559 -85
rect -497 85 -463 104
rect -497 17 -463 19
rect -497 -19 -463 -17
rect -497 -104 -463 -85
rect -401 85 -367 104
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -104 -367 -85
rect -305 85 -271 104
rect -305 17 -271 19
rect -305 -19 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 19
rect 271 -19 305 -17
rect 271 -104 305 -85
rect 367 85 401 104
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -104 401 -85
rect 463 85 497 104
rect 463 17 497 19
rect 463 -19 497 -17
rect 463 -104 497 -85
rect 559 85 593 104
rect 559 17 593 19
rect 559 -19 593 -17
rect 559 -104 593 -85
rect 655 85 689 104
rect 655 17 689 19
rect 655 -19 689 -17
rect 655 -104 689 -85
rect 751 85 785 104
rect 751 17 785 19
rect 751 -19 785 -17
rect 751 -104 785 -85
rect 847 85 881 104
rect 847 17 881 19
rect 847 -19 881 -17
rect 847 -104 881 -85
rect 943 85 977 104
rect 943 17 977 19
rect 943 -19 977 -17
rect 943 -104 977 -85
rect 1039 85 1073 104
rect 1039 17 1073 19
rect 1039 -19 1073 -17
rect 1039 -104 1073 -85
rect 1135 85 1169 104
rect 1135 17 1169 19
rect 1135 -19 1169 -17
rect 1135 -104 1169 -85
rect 1231 85 1265 104
rect 1231 17 1265 19
rect 1231 -19 1265 -17
rect 1231 -104 1265 -85
rect 1327 85 1361 104
rect 1327 17 1361 19
rect 1327 -19 1361 -17
rect 1327 -104 1361 -85
rect 1423 85 1457 104
rect 1423 17 1457 19
rect 1423 -19 1457 -17
rect 1423 -104 1457 -85
rect 1519 85 1553 104
rect 1519 17 1553 19
rect 1519 -19 1553 -17
rect 1519 -104 1553 -85
rect 1615 85 1649 104
rect 1615 17 1649 19
rect 1615 -19 1649 -17
rect 1615 -104 1649 -85
rect 1711 85 1745 104
rect 1711 17 1745 19
rect 1711 -19 1745 -17
rect 1711 -104 1745 -85
rect 1807 85 1841 104
rect 1807 17 1841 19
rect 1807 -19 1841 -17
rect 1807 -104 1841 -85
rect 1903 85 1937 104
rect 1903 17 1937 19
rect 1903 -19 1937 -17
rect 1903 -104 1937 -85
rect 1999 85 2033 104
rect 1999 17 2033 19
rect 1999 -19 2033 -17
rect 1999 -104 2033 -85
rect 2095 85 2129 104
rect 2095 17 2129 19
rect 2095 -19 2129 -17
rect 2095 -104 2129 -85
rect 2191 85 2225 104
rect 2191 17 2225 19
rect 2191 -19 2225 -17
rect 2191 -104 2225 -85
rect 2287 85 2321 104
rect 2287 17 2321 19
rect 2287 -19 2321 -17
rect 2287 -104 2321 -85
rect 2383 85 2417 104
rect 2383 17 2417 19
rect 2383 -19 2417 -17
rect 2383 -104 2417 -85
rect 2479 85 2513 104
rect 2479 17 2513 19
rect 2479 -19 2513 -17
rect 2479 -104 2513 -85
rect 2575 85 2609 104
rect 2575 17 2609 19
rect 2575 -19 2609 -17
rect 2575 -104 2609 -85
rect 2671 85 2705 104
rect 2671 17 2705 19
rect 2671 -19 2705 -17
rect 2671 -104 2705 -85
rect 2767 85 2801 104
rect 2767 17 2801 19
rect 2767 -19 2801 -17
rect 2767 -104 2801 -85
rect 2863 85 2897 104
rect 2863 17 2897 19
rect 2863 -19 2897 -17
rect 2863 -104 2897 -85
rect 2977 85 3011 119
rect 2977 17 3011 51
rect 2977 -51 3011 -17
rect 2977 -119 3011 -85
rect -3011 -240 -2977 -153
rect -2865 -172 -2849 -138
rect -2815 -172 -2799 -138
rect -2673 -172 -2657 -138
rect -2623 -172 -2607 -138
rect -2481 -172 -2465 -138
rect -2431 -172 -2415 -138
rect -2289 -172 -2273 -138
rect -2239 -172 -2223 -138
rect -2097 -172 -2081 -138
rect -2047 -172 -2031 -138
rect -1905 -172 -1889 -138
rect -1855 -172 -1839 -138
rect -1713 -172 -1697 -138
rect -1663 -172 -1647 -138
rect -1521 -172 -1505 -138
rect -1471 -172 -1455 -138
rect -1329 -172 -1313 -138
rect -1279 -172 -1263 -138
rect -1137 -172 -1121 -138
rect -1087 -172 -1071 -138
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 975 -172 991 -138
rect 1025 -172 1041 -138
rect 1167 -172 1183 -138
rect 1217 -172 1233 -138
rect 1359 -172 1375 -138
rect 1409 -172 1425 -138
rect 1551 -172 1567 -138
rect 1601 -172 1617 -138
rect 1743 -172 1759 -138
rect 1793 -172 1809 -138
rect 1935 -172 1951 -138
rect 1985 -172 2001 -138
rect 2127 -172 2143 -138
rect 2177 -172 2193 -138
rect 2319 -172 2335 -138
rect 2369 -172 2385 -138
rect 2511 -172 2527 -138
rect 2561 -172 2577 -138
rect 2703 -172 2719 -138
rect 2753 -172 2769 -138
rect 2977 -240 3011 -153
rect -3011 -274 -2907 -240
rect -2873 -274 -2839 -240
rect -2805 -274 -2771 -240
rect -2737 -274 -2703 -240
rect -2669 -274 -2635 -240
rect -2601 -274 -2567 -240
rect -2533 -274 -2499 -240
rect -2465 -274 -2431 -240
rect -2397 -274 -2363 -240
rect -2329 -274 -2295 -240
rect -2261 -274 -2227 -240
rect -2193 -274 -2159 -240
rect -2125 -274 -2091 -240
rect -2057 -274 -2023 -240
rect -1989 -274 -1955 -240
rect -1921 -274 -1887 -240
rect -1853 -274 -1819 -240
rect -1785 -274 -1751 -240
rect -1717 -274 -1683 -240
rect -1649 -274 -1615 -240
rect -1581 -274 -1547 -240
rect -1513 -274 -1479 -240
rect -1445 -274 -1411 -240
rect -1377 -274 -1343 -240
rect -1309 -274 -1275 -240
rect -1241 -274 -1207 -240
rect -1173 -274 -1139 -240
rect -1105 -274 -1071 -240
rect -1037 -274 -1003 -240
rect -969 -274 -935 -240
rect -901 -274 -867 -240
rect -833 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 833 -240
rect 867 -274 901 -240
rect 935 -274 969 -240
rect 1003 -274 1037 -240
rect 1071 -274 1105 -240
rect 1139 -274 1173 -240
rect 1207 -274 1241 -240
rect 1275 -274 1309 -240
rect 1343 -274 1377 -240
rect 1411 -274 1445 -240
rect 1479 -274 1513 -240
rect 1547 -274 1581 -240
rect 1615 -274 1649 -240
rect 1683 -274 1717 -240
rect 1751 -274 1785 -240
rect 1819 -274 1853 -240
rect 1887 -274 1921 -240
rect 1955 -274 1989 -240
rect 2023 -274 2057 -240
rect 2091 -274 2125 -240
rect 2159 -274 2193 -240
rect 2227 -274 2261 -240
rect 2295 -274 2329 -240
rect 2363 -274 2397 -240
rect 2431 -274 2465 -240
rect 2499 -274 2533 -240
rect 2567 -274 2601 -240
rect 2635 -274 2669 -240
rect 2703 -274 2737 -240
rect 2771 -274 2805 -240
rect 2839 -274 2873 -240
rect 2907 -274 3011 -240
<< viali >>
rect -2753 138 -2719 172
rect -2561 138 -2527 172
rect -2369 138 -2335 172
rect -2177 138 -2143 172
rect -1985 138 -1951 172
rect -1793 138 -1759 172
rect -1601 138 -1567 172
rect -1409 138 -1375 172
rect -1217 138 -1183 172
rect -1025 138 -991 172
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect 1087 138 1121 172
rect 1279 138 1313 172
rect 1471 138 1505 172
rect 1663 138 1697 172
rect 1855 138 1889 172
rect 2047 138 2081 172
rect 2239 138 2273 172
rect 2431 138 2465 172
rect 2623 138 2657 172
rect 2815 138 2849 172
rect -2897 51 -2863 53
rect -2897 19 -2863 51
rect -2897 -51 -2863 -19
rect -2897 -53 -2863 -51
rect -2801 51 -2767 53
rect -2801 19 -2767 51
rect -2801 -51 -2767 -19
rect -2801 -53 -2767 -51
rect -2705 51 -2671 53
rect -2705 19 -2671 51
rect -2705 -51 -2671 -19
rect -2705 -53 -2671 -51
rect -2609 51 -2575 53
rect -2609 19 -2575 51
rect -2609 -51 -2575 -19
rect -2609 -53 -2575 -51
rect -2513 51 -2479 53
rect -2513 19 -2479 51
rect -2513 -51 -2479 -19
rect -2513 -53 -2479 -51
rect -2417 51 -2383 53
rect -2417 19 -2383 51
rect -2417 -51 -2383 -19
rect -2417 -53 -2383 -51
rect -2321 51 -2287 53
rect -2321 19 -2287 51
rect -2321 -51 -2287 -19
rect -2321 -53 -2287 -51
rect -2225 51 -2191 53
rect -2225 19 -2191 51
rect -2225 -51 -2191 -19
rect -2225 -53 -2191 -51
rect -2129 51 -2095 53
rect -2129 19 -2095 51
rect -2129 -51 -2095 -19
rect -2129 -53 -2095 -51
rect -2033 51 -1999 53
rect -2033 19 -1999 51
rect -2033 -51 -1999 -19
rect -2033 -53 -1999 -51
rect -1937 51 -1903 53
rect -1937 19 -1903 51
rect -1937 -51 -1903 -19
rect -1937 -53 -1903 -51
rect -1841 51 -1807 53
rect -1841 19 -1807 51
rect -1841 -51 -1807 -19
rect -1841 -53 -1807 -51
rect -1745 51 -1711 53
rect -1745 19 -1711 51
rect -1745 -51 -1711 -19
rect -1745 -53 -1711 -51
rect -1649 51 -1615 53
rect -1649 19 -1615 51
rect -1649 -51 -1615 -19
rect -1649 -53 -1615 -51
rect -1553 51 -1519 53
rect -1553 19 -1519 51
rect -1553 -51 -1519 -19
rect -1553 -53 -1519 -51
rect -1457 51 -1423 53
rect -1457 19 -1423 51
rect -1457 -51 -1423 -19
rect -1457 -53 -1423 -51
rect -1361 51 -1327 53
rect -1361 19 -1327 51
rect -1361 -51 -1327 -19
rect -1361 -53 -1327 -51
rect -1265 51 -1231 53
rect -1265 19 -1231 51
rect -1265 -51 -1231 -19
rect -1265 -53 -1231 -51
rect -1169 51 -1135 53
rect -1169 19 -1135 51
rect -1169 -51 -1135 -19
rect -1169 -53 -1135 -51
rect -1073 51 -1039 53
rect -1073 19 -1039 51
rect -1073 -51 -1039 -19
rect -1073 -53 -1039 -51
rect -977 51 -943 53
rect -977 19 -943 51
rect -977 -51 -943 -19
rect -977 -53 -943 -51
rect -881 51 -847 53
rect -881 19 -847 51
rect -881 -51 -847 -19
rect -881 -53 -847 -51
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -689 51 -655 53
rect -689 19 -655 51
rect -689 -51 -655 -19
rect -689 -53 -655 -51
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 655 51 689 53
rect 655 19 689 51
rect 655 -51 689 -19
rect 655 -53 689 -51
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 847 51 881 53
rect 847 19 881 51
rect 847 -51 881 -19
rect 847 -53 881 -51
rect 943 51 977 53
rect 943 19 977 51
rect 943 -51 977 -19
rect 943 -53 977 -51
rect 1039 51 1073 53
rect 1039 19 1073 51
rect 1039 -51 1073 -19
rect 1039 -53 1073 -51
rect 1135 51 1169 53
rect 1135 19 1169 51
rect 1135 -51 1169 -19
rect 1135 -53 1169 -51
rect 1231 51 1265 53
rect 1231 19 1265 51
rect 1231 -51 1265 -19
rect 1231 -53 1265 -51
rect 1327 51 1361 53
rect 1327 19 1361 51
rect 1327 -51 1361 -19
rect 1327 -53 1361 -51
rect 1423 51 1457 53
rect 1423 19 1457 51
rect 1423 -51 1457 -19
rect 1423 -53 1457 -51
rect 1519 51 1553 53
rect 1519 19 1553 51
rect 1519 -51 1553 -19
rect 1519 -53 1553 -51
rect 1615 51 1649 53
rect 1615 19 1649 51
rect 1615 -51 1649 -19
rect 1615 -53 1649 -51
rect 1711 51 1745 53
rect 1711 19 1745 51
rect 1711 -51 1745 -19
rect 1711 -53 1745 -51
rect 1807 51 1841 53
rect 1807 19 1841 51
rect 1807 -51 1841 -19
rect 1807 -53 1841 -51
rect 1903 51 1937 53
rect 1903 19 1937 51
rect 1903 -51 1937 -19
rect 1903 -53 1937 -51
rect 1999 51 2033 53
rect 1999 19 2033 51
rect 1999 -51 2033 -19
rect 1999 -53 2033 -51
rect 2095 51 2129 53
rect 2095 19 2129 51
rect 2095 -51 2129 -19
rect 2095 -53 2129 -51
rect 2191 51 2225 53
rect 2191 19 2225 51
rect 2191 -51 2225 -19
rect 2191 -53 2225 -51
rect 2287 51 2321 53
rect 2287 19 2321 51
rect 2287 -51 2321 -19
rect 2287 -53 2321 -51
rect 2383 51 2417 53
rect 2383 19 2417 51
rect 2383 -51 2417 -19
rect 2383 -53 2417 -51
rect 2479 51 2513 53
rect 2479 19 2513 51
rect 2479 -51 2513 -19
rect 2479 -53 2513 -51
rect 2575 51 2609 53
rect 2575 19 2609 51
rect 2575 -51 2609 -19
rect 2575 -53 2609 -51
rect 2671 51 2705 53
rect 2671 19 2705 51
rect 2671 -51 2705 -19
rect 2671 -53 2705 -51
rect 2767 51 2801 53
rect 2767 19 2801 51
rect 2767 -51 2801 -19
rect 2767 -53 2801 -51
rect 2863 51 2897 53
rect 2863 19 2897 51
rect 2863 -51 2897 -19
rect 2863 -53 2897 -51
rect -2849 -172 -2815 -138
rect -2657 -172 -2623 -138
rect -2465 -172 -2431 -138
rect -2273 -172 -2239 -138
rect -2081 -172 -2047 -138
rect -1889 -172 -1855 -138
rect -1697 -172 -1663 -138
rect -1505 -172 -1471 -138
rect -1313 -172 -1279 -138
rect -1121 -172 -1087 -138
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
rect 991 -172 1025 -138
rect 1183 -172 1217 -138
rect 1375 -172 1409 -138
rect 1567 -172 1601 -138
rect 1759 -172 1793 -138
rect 1951 -172 1985 -138
rect 2143 -172 2177 -138
rect 2335 -172 2369 -138
rect 2527 -172 2561 -138
rect 2719 -172 2753 -138
<< metal1 >>
rect -2765 172 -2707 178
rect -2765 138 -2753 172
rect -2719 138 -2707 172
rect -2765 132 -2707 138
rect -2573 172 -2515 178
rect -2573 138 -2561 172
rect -2527 138 -2515 172
rect -2573 132 -2515 138
rect -2381 172 -2323 178
rect -2381 138 -2369 172
rect -2335 138 -2323 172
rect -2381 132 -2323 138
rect -2189 172 -2131 178
rect -2189 138 -2177 172
rect -2143 138 -2131 172
rect -2189 132 -2131 138
rect -1997 172 -1939 178
rect -1997 138 -1985 172
rect -1951 138 -1939 172
rect -1997 132 -1939 138
rect -1805 172 -1747 178
rect -1805 138 -1793 172
rect -1759 138 -1747 172
rect -1805 132 -1747 138
rect -1613 172 -1555 178
rect -1613 138 -1601 172
rect -1567 138 -1555 172
rect -1613 132 -1555 138
rect -1421 172 -1363 178
rect -1421 138 -1409 172
rect -1375 138 -1363 172
rect -1421 132 -1363 138
rect -1229 172 -1171 178
rect -1229 138 -1217 172
rect -1183 138 -1171 172
rect -1229 132 -1171 138
rect -1037 172 -979 178
rect -1037 138 -1025 172
rect -991 138 -979 172
rect -1037 132 -979 138
rect -845 172 -787 178
rect -845 138 -833 172
rect -799 138 -787 172
rect -845 132 -787 138
rect -653 172 -595 178
rect -653 138 -641 172
rect -607 138 -595 172
rect -653 132 -595 138
rect -461 172 -403 178
rect -461 138 -449 172
rect -415 138 -403 172
rect -461 132 -403 138
rect -269 172 -211 178
rect -269 138 -257 172
rect -223 138 -211 172
rect -269 132 -211 138
rect -77 172 -19 178
rect -77 138 -65 172
rect -31 138 -19 172
rect -77 132 -19 138
rect 115 172 173 178
rect 115 138 127 172
rect 161 138 173 172
rect 115 132 173 138
rect 307 172 365 178
rect 307 138 319 172
rect 353 138 365 172
rect 307 132 365 138
rect 499 172 557 178
rect 499 138 511 172
rect 545 138 557 172
rect 499 132 557 138
rect 691 172 749 178
rect 691 138 703 172
rect 737 138 749 172
rect 691 132 749 138
rect 883 172 941 178
rect 883 138 895 172
rect 929 138 941 172
rect 883 132 941 138
rect 1075 172 1133 178
rect 1075 138 1087 172
rect 1121 138 1133 172
rect 1075 132 1133 138
rect 1267 172 1325 178
rect 1267 138 1279 172
rect 1313 138 1325 172
rect 1267 132 1325 138
rect 1459 172 1517 178
rect 1459 138 1471 172
rect 1505 138 1517 172
rect 1459 132 1517 138
rect 1651 172 1709 178
rect 1651 138 1663 172
rect 1697 138 1709 172
rect 1651 132 1709 138
rect 1843 172 1901 178
rect 1843 138 1855 172
rect 1889 138 1901 172
rect 1843 132 1901 138
rect 2035 172 2093 178
rect 2035 138 2047 172
rect 2081 138 2093 172
rect 2035 132 2093 138
rect 2227 172 2285 178
rect 2227 138 2239 172
rect 2273 138 2285 172
rect 2227 132 2285 138
rect 2419 172 2477 178
rect 2419 138 2431 172
rect 2465 138 2477 172
rect 2419 132 2477 138
rect 2611 172 2669 178
rect 2611 138 2623 172
rect 2657 138 2669 172
rect 2611 132 2669 138
rect 2803 172 2861 178
rect 2803 138 2815 172
rect 2849 138 2861 172
rect 2803 132 2861 138
rect -2903 53 -2857 100
rect -2903 19 -2897 53
rect -2863 19 -2857 53
rect -2903 -19 -2857 19
rect -2903 -53 -2897 -19
rect -2863 -53 -2857 -19
rect -2903 -100 -2857 -53
rect -2807 53 -2761 100
rect -2807 19 -2801 53
rect -2767 19 -2761 53
rect -2807 -19 -2761 19
rect -2807 -53 -2801 -19
rect -2767 -53 -2761 -19
rect -2807 -100 -2761 -53
rect -2711 53 -2665 100
rect -2711 19 -2705 53
rect -2671 19 -2665 53
rect -2711 -19 -2665 19
rect -2711 -53 -2705 -19
rect -2671 -53 -2665 -19
rect -2711 -100 -2665 -53
rect -2615 53 -2569 100
rect -2615 19 -2609 53
rect -2575 19 -2569 53
rect -2615 -19 -2569 19
rect -2615 -53 -2609 -19
rect -2575 -53 -2569 -19
rect -2615 -100 -2569 -53
rect -2519 53 -2473 100
rect -2519 19 -2513 53
rect -2479 19 -2473 53
rect -2519 -19 -2473 19
rect -2519 -53 -2513 -19
rect -2479 -53 -2473 -19
rect -2519 -100 -2473 -53
rect -2423 53 -2377 100
rect -2423 19 -2417 53
rect -2383 19 -2377 53
rect -2423 -19 -2377 19
rect -2423 -53 -2417 -19
rect -2383 -53 -2377 -19
rect -2423 -100 -2377 -53
rect -2327 53 -2281 100
rect -2327 19 -2321 53
rect -2287 19 -2281 53
rect -2327 -19 -2281 19
rect -2327 -53 -2321 -19
rect -2287 -53 -2281 -19
rect -2327 -100 -2281 -53
rect -2231 53 -2185 100
rect -2231 19 -2225 53
rect -2191 19 -2185 53
rect -2231 -19 -2185 19
rect -2231 -53 -2225 -19
rect -2191 -53 -2185 -19
rect -2231 -100 -2185 -53
rect -2135 53 -2089 100
rect -2135 19 -2129 53
rect -2095 19 -2089 53
rect -2135 -19 -2089 19
rect -2135 -53 -2129 -19
rect -2095 -53 -2089 -19
rect -2135 -100 -2089 -53
rect -2039 53 -1993 100
rect -2039 19 -2033 53
rect -1999 19 -1993 53
rect -2039 -19 -1993 19
rect -2039 -53 -2033 -19
rect -1999 -53 -1993 -19
rect -2039 -100 -1993 -53
rect -1943 53 -1897 100
rect -1943 19 -1937 53
rect -1903 19 -1897 53
rect -1943 -19 -1897 19
rect -1943 -53 -1937 -19
rect -1903 -53 -1897 -19
rect -1943 -100 -1897 -53
rect -1847 53 -1801 100
rect -1847 19 -1841 53
rect -1807 19 -1801 53
rect -1847 -19 -1801 19
rect -1847 -53 -1841 -19
rect -1807 -53 -1801 -19
rect -1847 -100 -1801 -53
rect -1751 53 -1705 100
rect -1751 19 -1745 53
rect -1711 19 -1705 53
rect -1751 -19 -1705 19
rect -1751 -53 -1745 -19
rect -1711 -53 -1705 -19
rect -1751 -100 -1705 -53
rect -1655 53 -1609 100
rect -1655 19 -1649 53
rect -1615 19 -1609 53
rect -1655 -19 -1609 19
rect -1655 -53 -1649 -19
rect -1615 -53 -1609 -19
rect -1655 -100 -1609 -53
rect -1559 53 -1513 100
rect -1559 19 -1553 53
rect -1519 19 -1513 53
rect -1559 -19 -1513 19
rect -1559 -53 -1553 -19
rect -1519 -53 -1513 -19
rect -1559 -100 -1513 -53
rect -1463 53 -1417 100
rect -1463 19 -1457 53
rect -1423 19 -1417 53
rect -1463 -19 -1417 19
rect -1463 -53 -1457 -19
rect -1423 -53 -1417 -19
rect -1463 -100 -1417 -53
rect -1367 53 -1321 100
rect -1367 19 -1361 53
rect -1327 19 -1321 53
rect -1367 -19 -1321 19
rect -1367 -53 -1361 -19
rect -1327 -53 -1321 -19
rect -1367 -100 -1321 -53
rect -1271 53 -1225 100
rect -1271 19 -1265 53
rect -1231 19 -1225 53
rect -1271 -19 -1225 19
rect -1271 -53 -1265 -19
rect -1231 -53 -1225 -19
rect -1271 -100 -1225 -53
rect -1175 53 -1129 100
rect -1175 19 -1169 53
rect -1135 19 -1129 53
rect -1175 -19 -1129 19
rect -1175 -53 -1169 -19
rect -1135 -53 -1129 -19
rect -1175 -100 -1129 -53
rect -1079 53 -1033 100
rect -1079 19 -1073 53
rect -1039 19 -1033 53
rect -1079 -19 -1033 19
rect -1079 -53 -1073 -19
rect -1039 -53 -1033 -19
rect -1079 -100 -1033 -53
rect -983 53 -937 100
rect -983 19 -977 53
rect -943 19 -937 53
rect -983 -19 -937 19
rect -983 -53 -977 -19
rect -943 -53 -937 -19
rect -983 -100 -937 -53
rect -887 53 -841 100
rect -887 19 -881 53
rect -847 19 -841 53
rect -887 -19 -841 19
rect -887 -53 -881 -19
rect -847 -53 -841 -19
rect -887 -100 -841 -53
rect -791 53 -745 100
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -100 -745 -53
rect -695 53 -649 100
rect -695 19 -689 53
rect -655 19 -649 53
rect -695 -19 -649 19
rect -695 -53 -689 -19
rect -655 -53 -649 -19
rect -695 -100 -649 -53
rect -599 53 -553 100
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -100 -553 -53
rect -503 53 -457 100
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -100 -457 -53
rect -407 53 -361 100
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -100 -361 -53
rect -311 53 -265 100
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -100 -265 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 265 53 311 100
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -100 311 -53
rect 361 53 407 100
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -100 407 -53
rect 457 53 503 100
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -100 503 -53
rect 553 53 599 100
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -100 599 -53
rect 649 53 695 100
rect 649 19 655 53
rect 689 19 695 53
rect 649 -19 695 19
rect 649 -53 655 -19
rect 689 -53 695 -19
rect 649 -100 695 -53
rect 745 53 791 100
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -100 791 -53
rect 841 53 887 100
rect 841 19 847 53
rect 881 19 887 53
rect 841 -19 887 19
rect 841 -53 847 -19
rect 881 -53 887 -19
rect 841 -100 887 -53
rect 937 53 983 100
rect 937 19 943 53
rect 977 19 983 53
rect 937 -19 983 19
rect 937 -53 943 -19
rect 977 -53 983 -19
rect 937 -100 983 -53
rect 1033 53 1079 100
rect 1033 19 1039 53
rect 1073 19 1079 53
rect 1033 -19 1079 19
rect 1033 -53 1039 -19
rect 1073 -53 1079 -19
rect 1033 -100 1079 -53
rect 1129 53 1175 100
rect 1129 19 1135 53
rect 1169 19 1175 53
rect 1129 -19 1175 19
rect 1129 -53 1135 -19
rect 1169 -53 1175 -19
rect 1129 -100 1175 -53
rect 1225 53 1271 100
rect 1225 19 1231 53
rect 1265 19 1271 53
rect 1225 -19 1271 19
rect 1225 -53 1231 -19
rect 1265 -53 1271 -19
rect 1225 -100 1271 -53
rect 1321 53 1367 100
rect 1321 19 1327 53
rect 1361 19 1367 53
rect 1321 -19 1367 19
rect 1321 -53 1327 -19
rect 1361 -53 1367 -19
rect 1321 -100 1367 -53
rect 1417 53 1463 100
rect 1417 19 1423 53
rect 1457 19 1463 53
rect 1417 -19 1463 19
rect 1417 -53 1423 -19
rect 1457 -53 1463 -19
rect 1417 -100 1463 -53
rect 1513 53 1559 100
rect 1513 19 1519 53
rect 1553 19 1559 53
rect 1513 -19 1559 19
rect 1513 -53 1519 -19
rect 1553 -53 1559 -19
rect 1513 -100 1559 -53
rect 1609 53 1655 100
rect 1609 19 1615 53
rect 1649 19 1655 53
rect 1609 -19 1655 19
rect 1609 -53 1615 -19
rect 1649 -53 1655 -19
rect 1609 -100 1655 -53
rect 1705 53 1751 100
rect 1705 19 1711 53
rect 1745 19 1751 53
rect 1705 -19 1751 19
rect 1705 -53 1711 -19
rect 1745 -53 1751 -19
rect 1705 -100 1751 -53
rect 1801 53 1847 100
rect 1801 19 1807 53
rect 1841 19 1847 53
rect 1801 -19 1847 19
rect 1801 -53 1807 -19
rect 1841 -53 1847 -19
rect 1801 -100 1847 -53
rect 1897 53 1943 100
rect 1897 19 1903 53
rect 1937 19 1943 53
rect 1897 -19 1943 19
rect 1897 -53 1903 -19
rect 1937 -53 1943 -19
rect 1897 -100 1943 -53
rect 1993 53 2039 100
rect 1993 19 1999 53
rect 2033 19 2039 53
rect 1993 -19 2039 19
rect 1993 -53 1999 -19
rect 2033 -53 2039 -19
rect 1993 -100 2039 -53
rect 2089 53 2135 100
rect 2089 19 2095 53
rect 2129 19 2135 53
rect 2089 -19 2135 19
rect 2089 -53 2095 -19
rect 2129 -53 2135 -19
rect 2089 -100 2135 -53
rect 2185 53 2231 100
rect 2185 19 2191 53
rect 2225 19 2231 53
rect 2185 -19 2231 19
rect 2185 -53 2191 -19
rect 2225 -53 2231 -19
rect 2185 -100 2231 -53
rect 2281 53 2327 100
rect 2281 19 2287 53
rect 2321 19 2327 53
rect 2281 -19 2327 19
rect 2281 -53 2287 -19
rect 2321 -53 2327 -19
rect 2281 -100 2327 -53
rect 2377 53 2423 100
rect 2377 19 2383 53
rect 2417 19 2423 53
rect 2377 -19 2423 19
rect 2377 -53 2383 -19
rect 2417 -53 2423 -19
rect 2377 -100 2423 -53
rect 2473 53 2519 100
rect 2473 19 2479 53
rect 2513 19 2519 53
rect 2473 -19 2519 19
rect 2473 -53 2479 -19
rect 2513 -53 2519 -19
rect 2473 -100 2519 -53
rect 2569 53 2615 100
rect 2569 19 2575 53
rect 2609 19 2615 53
rect 2569 -19 2615 19
rect 2569 -53 2575 -19
rect 2609 -53 2615 -19
rect 2569 -100 2615 -53
rect 2665 53 2711 100
rect 2665 19 2671 53
rect 2705 19 2711 53
rect 2665 -19 2711 19
rect 2665 -53 2671 -19
rect 2705 -53 2711 -19
rect 2665 -100 2711 -53
rect 2761 53 2807 100
rect 2761 19 2767 53
rect 2801 19 2807 53
rect 2761 -19 2807 19
rect 2761 -53 2767 -19
rect 2801 -53 2807 -19
rect 2761 -100 2807 -53
rect 2857 53 2903 100
rect 2857 19 2863 53
rect 2897 19 2903 53
rect 2857 -19 2903 19
rect 2857 -53 2863 -19
rect 2897 -53 2903 -19
rect 2857 -100 2903 -53
rect -2861 -138 -2803 -132
rect -2861 -172 -2849 -138
rect -2815 -172 -2803 -138
rect -2861 -178 -2803 -172
rect -2669 -138 -2611 -132
rect -2669 -172 -2657 -138
rect -2623 -172 -2611 -138
rect -2669 -178 -2611 -172
rect -2477 -138 -2419 -132
rect -2477 -172 -2465 -138
rect -2431 -172 -2419 -138
rect -2477 -178 -2419 -172
rect -2285 -138 -2227 -132
rect -2285 -172 -2273 -138
rect -2239 -172 -2227 -138
rect -2285 -178 -2227 -172
rect -2093 -138 -2035 -132
rect -2093 -172 -2081 -138
rect -2047 -172 -2035 -138
rect -2093 -178 -2035 -172
rect -1901 -138 -1843 -132
rect -1901 -172 -1889 -138
rect -1855 -172 -1843 -138
rect -1901 -178 -1843 -172
rect -1709 -138 -1651 -132
rect -1709 -172 -1697 -138
rect -1663 -172 -1651 -138
rect -1709 -178 -1651 -172
rect -1517 -138 -1459 -132
rect -1517 -172 -1505 -138
rect -1471 -172 -1459 -138
rect -1517 -178 -1459 -172
rect -1325 -138 -1267 -132
rect -1325 -172 -1313 -138
rect -1279 -172 -1267 -138
rect -1325 -178 -1267 -172
rect -1133 -138 -1075 -132
rect -1133 -172 -1121 -138
rect -1087 -172 -1075 -138
rect -1133 -178 -1075 -172
rect -941 -138 -883 -132
rect -941 -172 -929 -138
rect -895 -172 -883 -138
rect -941 -178 -883 -172
rect -749 -138 -691 -132
rect -749 -172 -737 -138
rect -703 -172 -691 -138
rect -749 -178 -691 -172
rect -557 -138 -499 -132
rect -557 -172 -545 -138
rect -511 -172 -499 -138
rect -557 -178 -499 -172
rect -365 -138 -307 -132
rect -365 -172 -353 -138
rect -319 -172 -307 -138
rect -365 -178 -307 -172
rect -173 -138 -115 -132
rect -173 -172 -161 -138
rect -127 -172 -115 -138
rect -173 -178 -115 -172
rect 19 -138 77 -132
rect 19 -172 31 -138
rect 65 -172 77 -138
rect 19 -178 77 -172
rect 211 -138 269 -132
rect 211 -172 223 -138
rect 257 -172 269 -138
rect 211 -178 269 -172
rect 403 -138 461 -132
rect 403 -172 415 -138
rect 449 -172 461 -138
rect 403 -178 461 -172
rect 595 -138 653 -132
rect 595 -172 607 -138
rect 641 -172 653 -138
rect 595 -178 653 -172
rect 787 -138 845 -132
rect 787 -172 799 -138
rect 833 -172 845 -138
rect 787 -178 845 -172
rect 979 -138 1037 -132
rect 979 -172 991 -138
rect 1025 -172 1037 -138
rect 979 -178 1037 -172
rect 1171 -138 1229 -132
rect 1171 -172 1183 -138
rect 1217 -172 1229 -138
rect 1171 -178 1229 -172
rect 1363 -138 1421 -132
rect 1363 -172 1375 -138
rect 1409 -172 1421 -138
rect 1363 -178 1421 -172
rect 1555 -138 1613 -132
rect 1555 -172 1567 -138
rect 1601 -172 1613 -138
rect 1555 -178 1613 -172
rect 1747 -138 1805 -132
rect 1747 -172 1759 -138
rect 1793 -172 1805 -138
rect 1747 -178 1805 -172
rect 1939 -138 1997 -132
rect 1939 -172 1951 -138
rect 1985 -172 1997 -138
rect 1939 -178 1997 -172
rect 2131 -138 2189 -132
rect 2131 -172 2143 -138
rect 2177 -172 2189 -138
rect 2131 -178 2189 -172
rect 2323 -138 2381 -132
rect 2323 -172 2335 -138
rect 2369 -172 2381 -138
rect 2323 -178 2381 -172
rect 2515 -138 2573 -132
rect 2515 -172 2527 -138
rect 2561 -172 2573 -138
rect 2515 -178 2573 -172
rect 2707 -138 2765 -132
rect 2707 -172 2719 -138
rect 2753 -172 2765 -138
rect 2707 -178 2765 -172
<< properties >>
string FIXED_BBOX -2994 -257 2994 257
<< end >>
