magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -1117 -300 1117 300
<< nmoslvt >>
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
<< ndiff >>
rect -989 85 -927 100
rect -989 51 -977 85
rect -943 51 -927 85
rect -989 17 -927 51
rect -989 -17 -977 17
rect -943 -17 -927 17
rect -989 -51 -927 -17
rect -989 -85 -977 -51
rect -943 -85 -927 -51
rect -989 -100 -927 -85
rect -897 85 -831 100
rect -897 51 -881 85
rect -847 51 -831 85
rect -897 17 -831 51
rect -897 -17 -881 17
rect -847 -17 -831 17
rect -897 -51 -831 -17
rect -897 -85 -881 -51
rect -847 -85 -831 -51
rect -897 -100 -831 -85
rect -801 85 -735 100
rect -801 51 -785 85
rect -751 51 -735 85
rect -801 17 -735 51
rect -801 -17 -785 17
rect -751 -17 -735 17
rect -801 -51 -735 -17
rect -801 -85 -785 -51
rect -751 -85 -735 -51
rect -801 -100 -735 -85
rect -705 85 -639 100
rect -705 51 -689 85
rect -655 51 -639 85
rect -705 17 -639 51
rect -705 -17 -689 17
rect -655 -17 -639 17
rect -705 -51 -639 -17
rect -705 -85 -689 -51
rect -655 -85 -639 -51
rect -705 -100 -639 -85
rect -609 85 -543 100
rect -609 51 -593 85
rect -559 51 -543 85
rect -609 17 -543 51
rect -609 -17 -593 17
rect -559 -17 -543 17
rect -609 -51 -543 -17
rect -609 -85 -593 -51
rect -559 -85 -543 -51
rect -609 -100 -543 -85
rect -513 85 -447 100
rect -513 51 -497 85
rect -463 51 -447 85
rect -513 17 -447 51
rect -513 -17 -497 17
rect -463 -17 -447 17
rect -513 -51 -447 -17
rect -513 -85 -497 -51
rect -463 -85 -447 -51
rect -513 -100 -447 -85
rect -417 85 -351 100
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -100 -351 -85
rect -321 85 -255 100
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 321 100
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -100 321 -85
rect 351 85 417 100
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -100 417 -85
rect 447 85 513 100
rect 447 51 463 85
rect 497 51 513 85
rect 447 17 513 51
rect 447 -17 463 17
rect 497 -17 513 17
rect 447 -51 513 -17
rect 447 -85 463 -51
rect 497 -85 513 -51
rect 447 -100 513 -85
rect 543 85 609 100
rect 543 51 559 85
rect 593 51 609 85
rect 543 17 609 51
rect 543 -17 559 17
rect 593 -17 609 17
rect 543 -51 609 -17
rect 543 -85 559 -51
rect 593 -85 609 -51
rect 543 -100 609 -85
rect 639 85 705 100
rect 639 51 655 85
rect 689 51 705 85
rect 639 17 705 51
rect 639 -17 655 17
rect 689 -17 705 17
rect 639 -51 705 -17
rect 639 -85 655 -51
rect 689 -85 705 -51
rect 639 -100 705 -85
rect 735 85 801 100
rect 735 51 751 85
rect 785 51 801 85
rect 735 17 801 51
rect 735 -17 751 17
rect 785 -17 801 17
rect 735 -51 801 -17
rect 735 -85 751 -51
rect 785 -85 801 -51
rect 735 -100 801 -85
rect 831 85 897 100
rect 831 51 847 85
rect 881 51 897 85
rect 831 17 897 51
rect 831 -17 847 17
rect 881 -17 897 17
rect 831 -51 897 -17
rect 831 -85 847 -51
rect 881 -85 897 -51
rect 831 -100 897 -85
rect 927 85 989 100
rect 927 51 943 85
rect 977 51 989 85
rect 927 17 989 51
rect 927 -17 943 17
rect 977 -17 989 17
rect 927 -51 989 -17
rect 927 -85 943 -51
rect 977 -85 989 -51
rect 927 -100 989 -85
<< ndiffc >>
rect -977 51 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -51
rect -881 51 -847 85
rect -881 -17 -847 17
rect -881 -85 -847 -51
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -689 51 -655 85
rect -689 -17 -655 17
rect -689 -85 -655 -51
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 655 51 689 85
rect 655 -17 689 17
rect 655 -85 689 -51
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 847 51 881 85
rect 847 -17 881 17
rect 847 -85 881 -51
rect 943 51 977 85
rect 943 -17 977 17
rect 943 -85 977 -51
<< psubdiff >>
rect -1091 240 -969 274
rect -935 240 -901 274
rect -867 240 -833 274
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect 833 240 867 274
rect 901 240 935 274
rect 969 240 1091 274
rect -1091 153 -1057 240
rect -1091 85 -1057 119
rect 1057 153 1091 240
rect -1091 17 -1057 51
rect -1091 -51 -1057 -17
rect -1091 -119 -1057 -85
rect 1057 85 1091 119
rect 1057 17 1091 51
rect 1057 -51 1091 -17
rect -1091 -240 -1057 -153
rect 1057 -119 1091 -85
rect 1057 -240 1091 -153
rect -1091 -274 -969 -240
rect -935 -274 -901 -240
rect -867 -274 -833 -240
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
rect 833 -274 867 -240
rect 901 -274 935 -240
rect 969 -274 1091 -240
<< psubdiffcont >>
rect -969 240 -935 274
rect -901 240 -867 274
rect -833 240 -799 274
rect -765 240 -731 274
rect -697 240 -663 274
rect -629 240 -595 274
rect -561 240 -527 274
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect 527 240 561 274
rect 595 240 629 274
rect 663 240 697 274
rect 731 240 765 274
rect 799 240 833 274
rect 867 240 901 274
rect 935 240 969 274
rect -1091 119 -1057 153
rect 1057 119 1091 153
rect -1091 51 -1057 85
rect -1091 -17 -1057 17
rect -1091 -85 -1057 -51
rect 1057 51 1091 85
rect 1057 -17 1091 17
rect 1057 -85 1091 -51
rect -1091 -153 -1057 -119
rect 1057 -153 1091 -119
rect -969 -274 -935 -240
rect -901 -274 -867 -240
rect -833 -274 -799 -240
rect -765 -274 -731 -240
rect -697 -274 -663 -240
rect -629 -274 -595 -240
rect -561 -274 -527 -240
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
rect 527 -274 561 -240
rect 595 -274 629 -240
rect 663 -274 697 -240
rect 731 -274 765 -240
rect 799 -274 833 -240
rect 867 -274 901 -240
rect 935 -274 969 -240
<< poly >>
rect -849 172 -783 188
rect -849 138 -833 172
rect -799 138 -783 172
rect -927 100 -897 126
rect -849 122 -783 138
rect -657 172 -591 188
rect -657 138 -641 172
rect -607 138 -591 172
rect -831 100 -801 122
rect -735 100 -705 126
rect -657 122 -591 138
rect -465 172 -399 188
rect -465 138 -449 172
rect -415 138 -399 172
rect -639 100 -609 122
rect -543 100 -513 126
rect -465 122 -399 138
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -447 100 -417 122
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 495 172 561 188
rect 495 138 511 172
rect 545 138 561 172
rect 321 100 351 122
rect 417 100 447 126
rect 495 122 561 138
rect 687 172 753 188
rect 687 138 703 172
rect 737 138 753 172
rect 513 100 543 122
rect 609 100 639 126
rect 687 122 753 138
rect 879 172 945 188
rect 879 138 895 172
rect 929 138 945 172
rect 705 100 735 122
rect 801 100 831 126
rect 879 122 945 138
rect 897 100 927 122
rect -927 -122 -897 -100
rect -945 -138 -879 -122
rect -831 -126 -801 -100
rect -735 -122 -705 -100
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -945 -188 -879 -172
rect -753 -138 -687 -122
rect -639 -126 -609 -100
rect -543 -122 -513 -100
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -753 -188 -687 -172
rect -561 -138 -495 -122
rect -447 -126 -417 -100
rect -351 -122 -321 -100
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -561 -188 -495 -172
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 417 -122 447 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
rect 399 -138 465 -122
rect 513 -126 543 -100
rect 609 -122 639 -100
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 399 -188 465 -172
rect 591 -138 657 -122
rect 705 -126 735 -100
rect 801 -122 831 -100
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 591 -188 657 -172
rect 783 -138 849 -122
rect 897 -126 927 -100
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 783 -188 849 -172
<< polycont >>
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
<< locali >>
rect -1091 240 -969 274
rect -935 240 -901 274
rect -867 240 -833 274
rect -799 240 -765 274
rect -731 240 -697 274
rect -663 240 -629 274
rect -595 240 -561 274
rect -527 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 527 274
rect 561 240 595 274
rect 629 240 663 274
rect 697 240 731 274
rect 765 240 799 274
rect 833 240 867 274
rect 901 240 935 274
rect 969 240 1091 274
rect -1091 153 -1057 240
rect -849 138 -833 172
rect -799 138 -783 172
rect -657 138 -641 172
rect -607 138 -591 172
rect -465 138 -449 172
rect -415 138 -399 172
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect 495 138 511 172
rect 545 138 561 172
rect 687 138 703 172
rect 737 138 753 172
rect 879 138 895 172
rect 929 138 945 172
rect 1057 153 1091 240
rect -1091 85 -1057 119
rect -1091 17 -1057 51
rect -1091 -51 -1057 -17
rect -1091 -119 -1057 -85
rect -977 85 -943 104
rect -977 17 -943 19
rect -977 -19 -943 -17
rect -977 -104 -943 -85
rect -881 85 -847 104
rect -881 17 -847 19
rect -881 -19 -847 -17
rect -881 -104 -847 -85
rect -785 85 -751 104
rect -785 17 -751 19
rect -785 -19 -751 -17
rect -785 -104 -751 -85
rect -689 85 -655 104
rect -689 17 -655 19
rect -689 -19 -655 -17
rect -689 -104 -655 -85
rect -593 85 -559 104
rect -593 17 -559 19
rect -593 -19 -559 -17
rect -593 -104 -559 -85
rect -497 85 -463 104
rect -497 17 -463 19
rect -497 -19 -463 -17
rect -497 -104 -463 -85
rect -401 85 -367 104
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -104 -367 -85
rect -305 85 -271 104
rect -305 17 -271 19
rect -305 -19 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 19
rect 271 -19 305 -17
rect 271 -104 305 -85
rect 367 85 401 104
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -104 401 -85
rect 463 85 497 104
rect 463 17 497 19
rect 463 -19 497 -17
rect 463 -104 497 -85
rect 559 85 593 104
rect 559 17 593 19
rect 559 -19 593 -17
rect 559 -104 593 -85
rect 655 85 689 104
rect 655 17 689 19
rect 655 -19 689 -17
rect 655 -104 689 -85
rect 751 85 785 104
rect 751 17 785 19
rect 751 -19 785 -17
rect 751 -104 785 -85
rect 847 85 881 104
rect 847 17 881 19
rect 847 -19 881 -17
rect 847 -104 881 -85
rect 943 85 977 104
rect 943 17 977 19
rect 943 -19 977 -17
rect 943 -104 977 -85
rect 1057 85 1091 119
rect 1057 17 1091 51
rect 1057 -51 1091 -17
rect 1057 -119 1091 -85
rect -1091 -240 -1057 -153
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 1057 -240 1091 -153
rect -1091 -274 -969 -240
rect -935 -274 -901 -240
rect -867 -274 -833 -240
rect -799 -274 -765 -240
rect -731 -274 -697 -240
rect -663 -274 -629 -240
rect -595 -274 -561 -240
rect -527 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 527 -240
rect 561 -274 595 -240
rect 629 -274 663 -240
rect 697 -274 731 -240
rect 765 -274 799 -240
rect 833 -274 867 -240
rect 901 -274 935 -240
rect 969 -274 1091 -240
<< viali >>
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect -977 51 -943 53
rect -977 19 -943 51
rect -977 -51 -943 -19
rect -977 -53 -943 -51
rect -881 51 -847 53
rect -881 19 -847 51
rect -881 -51 -847 -19
rect -881 -53 -847 -51
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -689 51 -655 53
rect -689 19 -655 51
rect -689 -51 -655 -19
rect -689 -53 -655 -51
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 655 51 689 53
rect 655 19 689 51
rect 655 -51 689 -19
rect 655 -53 689 -51
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 847 51 881 53
rect 847 19 881 51
rect 847 -51 881 -19
rect 847 -53 881 -51
rect 943 51 977 53
rect 943 19 977 51
rect 943 -51 977 -19
rect 943 -53 977 -51
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
<< metal1 >>
rect -845 175 -787 178
rect -653 175 -595 178
rect -461 175 -403 178
rect -269 175 -211 178
rect -77 175 -19 178
rect 115 175 173 178
rect 307 175 365 178
rect 499 175 557 178
rect 691 175 749 178
rect 883 175 941 178
rect -850 172 1090 175
rect -850 140 -833 172
rect -845 138 -833 140
rect -799 140 -641 172
rect -799 138 -787 140
rect -845 132 -787 138
rect -653 138 -641 140
rect -607 140 -449 172
rect -607 138 -595 140
rect -653 132 -595 138
rect -461 138 -449 140
rect -415 140 -257 172
rect -415 138 -403 140
rect -461 132 -403 138
rect -269 138 -257 140
rect -223 140 -65 172
rect -223 138 -211 140
rect -269 132 -211 138
rect -77 138 -65 140
rect -31 140 127 172
rect -31 138 -19 140
rect -77 132 -19 138
rect 115 138 127 140
rect 161 140 319 172
rect 161 138 173 140
rect 115 132 173 138
rect 307 138 319 140
rect 353 140 511 172
rect 353 138 365 140
rect 307 132 365 138
rect 499 138 511 140
rect 545 140 703 172
rect 545 138 557 140
rect 499 132 557 138
rect 691 138 703 140
rect 737 140 895 172
rect 737 138 749 140
rect 691 132 749 138
rect 883 138 895 140
rect 929 140 1090 172
rect 929 138 941 140
rect 883 132 941 138
rect -983 53 -937 100
rect -983 19 -977 53
rect -943 19 -937 53
rect -983 -19 -937 19
rect -983 -53 -977 -19
rect -943 -53 -937 -19
rect -983 -100 -937 -53
rect -887 53 -841 100
rect -887 19 -881 53
rect -847 19 -841 53
rect -887 -19 -841 19
rect -887 -53 -881 -19
rect -847 -53 -841 -19
rect -887 -100 -841 -53
rect -791 53 -745 100
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -100 -745 -53
rect -695 53 -649 100
rect -695 19 -689 53
rect -655 19 -649 53
rect -695 -19 -649 19
rect -695 -53 -689 -19
rect -655 -53 -649 -19
rect -695 -100 -649 -53
rect -599 53 -553 100
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -100 -553 -53
rect -503 53 -457 100
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -100 -457 -53
rect -407 53 -361 100
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -100 -361 -53
rect -311 53 -265 100
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -100 -265 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 265 53 311 100
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -100 311 -53
rect 361 53 407 100
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -100 407 -53
rect 457 53 503 100
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -100 503 -53
rect 553 53 599 100
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -100 599 -53
rect 649 53 695 100
rect 649 19 655 53
rect 689 19 695 53
rect 649 -19 695 19
rect 649 -53 655 -19
rect 689 -53 695 -19
rect 649 -100 695 -53
rect 745 53 791 100
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -100 791 -53
rect 841 53 887 100
rect 841 19 847 53
rect 881 19 887 53
rect 841 -19 887 19
rect 841 -53 847 -19
rect 881 -53 887 -19
rect 841 -100 887 -53
rect 937 53 983 100
rect 937 19 943 53
rect 977 19 983 53
rect 937 -19 983 19
rect 937 -53 943 -19
rect 977 -53 983 -19
rect 937 -100 983 -53
rect -941 -138 -883 -132
rect -941 -140 -929 -138
rect -945 -172 -929 -140
rect -895 -140 -883 -138
rect -749 -138 -691 -132
rect -749 -140 -737 -138
rect -895 -172 -737 -140
rect -703 -140 -691 -138
rect -557 -138 -499 -132
rect -557 -140 -545 -138
rect -703 -172 -545 -140
rect -511 -140 -499 -138
rect -365 -138 -307 -132
rect -365 -140 -353 -138
rect -511 -172 -353 -140
rect -319 -140 -307 -138
rect -173 -138 -115 -132
rect -173 -140 -161 -138
rect -319 -172 -161 -140
rect -127 -140 -115 -138
rect 19 -138 77 -132
rect 19 -140 31 -138
rect -127 -172 31 -140
rect 65 -140 77 -138
rect 211 -138 269 -132
rect 211 -140 223 -138
rect 65 -172 223 -140
rect 257 -140 269 -138
rect 403 -138 461 -132
rect 403 -140 415 -138
rect 257 -172 415 -140
rect 449 -140 461 -138
rect 595 -138 653 -132
rect 595 -140 607 -138
rect 449 -172 607 -140
rect 641 -140 653 -138
rect 787 -138 845 -132
rect 787 -140 799 -138
rect 641 -172 799 -140
rect 833 -140 845 -138
rect 1060 -140 1090 140
rect 833 -172 1090 -140
rect -945 -175 1090 -172
rect -941 -178 -883 -175
rect -749 -178 -691 -175
rect -557 -178 -499 -175
rect -365 -178 -307 -175
rect -173 -178 -115 -175
rect 19 -178 77 -175
rect 211 -178 269 -175
rect 403 -178 461 -175
rect 595 -178 653 -175
rect 787 -178 845 -175
<< properties >>
string FIXED_BBOX -1074 -257 1074 257
<< end >>
