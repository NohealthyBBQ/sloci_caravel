magic
tech sky130A
timestamp 1669931839
<< locali >>
rect -11930 -65060 -11680 -65040
rect -11930 -65190 -11680 -65170
rect -11930 -65320 -11680 -65300
<< metal1 >>
rect -12000 7500 110000 12000
rect -12000 4500 500 7500
rect 99500 4500 110000 7500
rect -12000 -1500 110000 4500
rect -12000 -4500 500 -1500
rect 99500 -4500 110000 -1500
rect -12000 -9000 110000 -4500
rect -12000 -39000 0 -9000
rect 100000 -39000 110000 -9000
rect -12000 -54500 110000 -39000
rect -12000 -57500 500 -54500
rect 99500 -57500 110000 -54500
rect -12000 -64000 110000 -57500
<< via1 >>
rect 500 4500 99500 7500
rect 500 -4500 99500 -1500
rect 500 -57500 99500 -54500
<< metal2 >>
rect 0 7500 100000 8000
rect 0 4500 500 7500
rect 99500 4500 100000 7500
rect 0 4000 100000 4500
rect 0 -1500 100000 -1000
rect 0 -4500 500 -1500
rect 99500 -4500 100000 -1500
rect 0 -5000 100000 -4500
rect 0 -45500 100000 -45000
rect 0 -48500 500 -45500
rect 99500 -48500 100000 -45500
rect 0 -49000 100000 -48500
rect 0 -54500 100000 -54000
rect 0 -57500 500 -54500
rect 99500 -57500 100000 -54500
rect 0 -58000 100000 -57500
<< via2 >>
rect 500 4500 99500 7500
rect 500 -4500 99500 -1500
rect 500 -48500 99500 -45500
rect 500 -57500 99500 -54500
<< metal3 >>
rect 0 7500 100000 8000
rect 0 4500 500 7500
rect 99500 4500 100000 7500
rect 0 4000 100000 4500
rect 0 -1500 100000 -1000
rect 0 -4500 500 -1500
rect 99500 -4500 100000 -1500
rect 0 -5000 100000 -4500
rect 0 -45500 100000 -45000
rect 0 -48500 500 -45500
rect 99500 -48500 100000 -45500
rect 0 -49000 100000 -48500
rect 0 -54500 100000 -54000
rect 0 -57500 500 -54500
rect 99500 -57500 100000 -54500
rect 0 -58000 100000 -57500
<< via3 >>
rect 500 4500 99500 7500
rect 500 -4500 99500 -1500
rect 500 -48500 99500 -45500
rect 500 -57500 99500 -54500
<< metal4 >>
rect 0 7500 100000 8000
rect 0 4500 500 7500
rect 99500 4500 100000 7500
rect 0 4000 100000 4500
rect 0 -1500 100000 -1000
rect 0 -4500 500 -1500
rect 99500 -4500 100000 -1500
rect 0 -5000 100000 -4500
rect 0 -45500 100000 -45000
rect 0 -48500 500 -45500
rect 99500 -48500 100000 -45500
rect 0 -49000 100000 -48500
rect 0 -54500 100000 -54000
rect 0 -57500 500 -54500
rect 99500 -57500 100000 -54500
rect 0 -58000 100000 -57500
<< via4 >>
rect 500 4500 99500 7500
rect 500 -4500 99500 -1500
rect 500 -48500 99500 -45500
rect 500 -57500 99500 -54500
<< metal5 >>
rect 0 7500 100000 8000
rect 0 4500 500 7500
rect 99500 4500 100000 7500
rect 0 4000 100000 4500
rect -1000 1000 101000 2000
rect 0 -1500 100000 -1000
rect 0 -4500 500 -1500
rect 99500 -4500 100000 -1500
rect 0 -5000 100000 -4500
rect 0 -45500 100000 -45000
rect 0 -48500 500 -45500
rect 99500 -48500 100000 -45500
rect 0 -49000 100000 -48500
rect -1000 -52000 100000 -51000
rect 0 -54500 100000 -54000
rect 0 -57500 500 -54500
rect 99500 -57500 100000 -54500
rect 0 -58000 100000 -57500
use sky130_fd_pr__nfet_01v8_lvt_M9466H  sky130_fd_pr__nfet_01v8_lvt_M9466H_0
timestamp 1669931839
transform 1 0 -11805 0 1 -65180
box -148 -205 148 205
<< labels >>
flabel metal1 -12000 -64000 110000 -57500 0 FreeSans 20000 0 0 0 GND
flabel metal5 -1000 1000 0 2000 0 FreeSans 20000 0 0 0 INA
flabel metal5 100000 1000 101000 2000 0 FreeSans 20000 0 0 0 OUTA
flabel metal5 -1000 -52000 0 -51000 0 FreeSans 20000 0 0 0 INB
flabel metal1 100000 -52000 101000 -51000 0 FreeSans 20000 0 0 0 OUTB
<< end >>
