magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -441 4702 441 4788
rect -441 -4702 -355 4702
rect 355 -4702 441 4702
rect -441 -4788 441 -4702
<< psubdiff >>
rect -415 4728 -289 4762
rect -255 4728 -221 4762
rect -187 4728 -153 4762
rect -119 4728 -85 4762
rect -51 4728 -17 4762
rect 17 4728 51 4762
rect 85 4728 119 4762
rect 153 4728 187 4762
rect 221 4728 255 4762
rect 289 4728 415 4762
rect -415 4641 -381 4728
rect 381 4641 415 4728
rect -415 4573 -381 4607
rect -415 4505 -381 4539
rect -415 4437 -381 4471
rect -415 4369 -381 4403
rect -415 4301 -381 4335
rect -415 4233 -381 4267
rect -415 4165 -381 4199
rect -415 4097 -381 4131
rect -415 4029 -381 4063
rect -415 3961 -381 3995
rect -415 3893 -381 3927
rect -415 3825 -381 3859
rect -415 3757 -381 3791
rect -415 3689 -381 3723
rect -415 3621 -381 3655
rect -415 3553 -381 3587
rect -415 3485 -381 3519
rect -415 3417 -381 3451
rect -415 3349 -381 3383
rect -415 3281 -381 3315
rect -415 3213 -381 3247
rect -415 3145 -381 3179
rect -415 3077 -381 3111
rect -415 3009 -381 3043
rect -415 2941 -381 2975
rect -415 2873 -381 2907
rect -415 2805 -381 2839
rect -415 2737 -381 2771
rect -415 2669 -381 2703
rect -415 2601 -381 2635
rect -415 2533 -381 2567
rect -415 2465 -381 2499
rect -415 2397 -381 2431
rect -415 2329 -381 2363
rect -415 2261 -381 2295
rect -415 2193 -381 2227
rect -415 2125 -381 2159
rect -415 2057 -381 2091
rect -415 1989 -381 2023
rect -415 1921 -381 1955
rect -415 1853 -381 1887
rect -415 1785 -381 1819
rect -415 1717 -381 1751
rect -415 1649 -381 1683
rect -415 1581 -381 1615
rect -415 1513 -381 1547
rect -415 1445 -381 1479
rect -415 1377 -381 1411
rect -415 1309 -381 1343
rect -415 1241 -381 1275
rect -415 1173 -381 1207
rect -415 1105 -381 1139
rect -415 1037 -381 1071
rect -415 969 -381 1003
rect -415 901 -381 935
rect -415 833 -381 867
rect -415 765 -381 799
rect -415 697 -381 731
rect -415 629 -381 663
rect -415 561 -381 595
rect -415 493 -381 527
rect -415 425 -381 459
rect -415 357 -381 391
rect -415 289 -381 323
rect -415 221 -381 255
rect -415 153 -381 187
rect -415 85 -381 119
rect -415 17 -381 51
rect -415 -51 -381 -17
rect -415 -119 -381 -85
rect -415 -187 -381 -153
rect -415 -255 -381 -221
rect -415 -323 -381 -289
rect -415 -391 -381 -357
rect -415 -459 -381 -425
rect -415 -527 -381 -493
rect -415 -595 -381 -561
rect -415 -663 -381 -629
rect -415 -731 -381 -697
rect -415 -799 -381 -765
rect -415 -867 -381 -833
rect -415 -935 -381 -901
rect -415 -1003 -381 -969
rect -415 -1071 -381 -1037
rect -415 -1139 -381 -1105
rect -415 -1207 -381 -1173
rect -415 -1275 -381 -1241
rect -415 -1343 -381 -1309
rect -415 -1411 -381 -1377
rect -415 -1479 -381 -1445
rect -415 -1547 -381 -1513
rect -415 -1615 -381 -1581
rect -415 -1683 -381 -1649
rect -415 -1751 -381 -1717
rect -415 -1819 -381 -1785
rect -415 -1887 -381 -1853
rect -415 -1955 -381 -1921
rect -415 -2023 -381 -1989
rect -415 -2091 -381 -2057
rect -415 -2159 -381 -2125
rect -415 -2227 -381 -2193
rect -415 -2295 -381 -2261
rect -415 -2363 -381 -2329
rect -415 -2431 -381 -2397
rect -415 -2499 -381 -2465
rect -415 -2567 -381 -2533
rect -415 -2635 -381 -2601
rect -415 -2703 -381 -2669
rect -415 -2771 -381 -2737
rect -415 -2839 -381 -2805
rect -415 -2907 -381 -2873
rect -415 -2975 -381 -2941
rect -415 -3043 -381 -3009
rect -415 -3111 -381 -3077
rect -415 -3179 -381 -3145
rect -415 -3247 -381 -3213
rect -415 -3315 -381 -3281
rect -415 -3383 -381 -3349
rect -415 -3451 -381 -3417
rect -415 -3519 -381 -3485
rect -415 -3587 -381 -3553
rect -415 -3655 -381 -3621
rect -415 -3723 -381 -3689
rect -415 -3791 -381 -3757
rect -415 -3859 -381 -3825
rect -415 -3927 -381 -3893
rect -415 -3995 -381 -3961
rect -415 -4063 -381 -4029
rect -415 -4131 -381 -4097
rect -415 -4199 -381 -4165
rect -415 -4267 -381 -4233
rect -415 -4335 -381 -4301
rect -415 -4403 -381 -4369
rect -415 -4471 -381 -4437
rect -415 -4539 -381 -4505
rect -415 -4607 -381 -4573
rect 381 4573 415 4607
rect 381 4505 415 4539
rect 381 4437 415 4471
rect 381 4369 415 4403
rect 381 4301 415 4335
rect 381 4233 415 4267
rect 381 4165 415 4199
rect 381 4097 415 4131
rect 381 4029 415 4063
rect 381 3961 415 3995
rect 381 3893 415 3927
rect 381 3825 415 3859
rect 381 3757 415 3791
rect 381 3689 415 3723
rect 381 3621 415 3655
rect 381 3553 415 3587
rect 381 3485 415 3519
rect 381 3417 415 3451
rect 381 3349 415 3383
rect 381 3281 415 3315
rect 381 3213 415 3247
rect 381 3145 415 3179
rect 381 3077 415 3111
rect 381 3009 415 3043
rect 381 2941 415 2975
rect 381 2873 415 2907
rect 381 2805 415 2839
rect 381 2737 415 2771
rect 381 2669 415 2703
rect 381 2601 415 2635
rect 381 2533 415 2567
rect 381 2465 415 2499
rect 381 2397 415 2431
rect 381 2329 415 2363
rect 381 2261 415 2295
rect 381 2193 415 2227
rect 381 2125 415 2159
rect 381 2057 415 2091
rect 381 1989 415 2023
rect 381 1921 415 1955
rect 381 1853 415 1887
rect 381 1785 415 1819
rect 381 1717 415 1751
rect 381 1649 415 1683
rect 381 1581 415 1615
rect 381 1513 415 1547
rect 381 1445 415 1479
rect 381 1377 415 1411
rect 381 1309 415 1343
rect 381 1241 415 1275
rect 381 1173 415 1207
rect 381 1105 415 1139
rect 381 1037 415 1071
rect 381 969 415 1003
rect 381 901 415 935
rect 381 833 415 867
rect 381 765 415 799
rect 381 697 415 731
rect 381 629 415 663
rect 381 561 415 595
rect 381 493 415 527
rect 381 425 415 459
rect 381 357 415 391
rect 381 289 415 323
rect 381 221 415 255
rect 381 153 415 187
rect 381 85 415 119
rect 381 17 415 51
rect 381 -51 415 -17
rect 381 -119 415 -85
rect 381 -187 415 -153
rect 381 -255 415 -221
rect 381 -323 415 -289
rect 381 -391 415 -357
rect 381 -459 415 -425
rect 381 -527 415 -493
rect 381 -595 415 -561
rect 381 -663 415 -629
rect 381 -731 415 -697
rect 381 -799 415 -765
rect 381 -867 415 -833
rect 381 -935 415 -901
rect 381 -1003 415 -969
rect 381 -1071 415 -1037
rect 381 -1139 415 -1105
rect 381 -1207 415 -1173
rect 381 -1275 415 -1241
rect 381 -1343 415 -1309
rect 381 -1411 415 -1377
rect 381 -1479 415 -1445
rect 381 -1547 415 -1513
rect 381 -1615 415 -1581
rect 381 -1683 415 -1649
rect 381 -1751 415 -1717
rect 381 -1819 415 -1785
rect 381 -1887 415 -1853
rect 381 -1955 415 -1921
rect 381 -2023 415 -1989
rect 381 -2091 415 -2057
rect 381 -2159 415 -2125
rect 381 -2227 415 -2193
rect 381 -2295 415 -2261
rect 381 -2363 415 -2329
rect 381 -2431 415 -2397
rect 381 -2499 415 -2465
rect 381 -2567 415 -2533
rect 381 -2635 415 -2601
rect 381 -2703 415 -2669
rect 381 -2771 415 -2737
rect 381 -2839 415 -2805
rect 381 -2907 415 -2873
rect 381 -2975 415 -2941
rect 381 -3043 415 -3009
rect 381 -3111 415 -3077
rect 381 -3179 415 -3145
rect 381 -3247 415 -3213
rect 381 -3315 415 -3281
rect 381 -3383 415 -3349
rect 381 -3451 415 -3417
rect 381 -3519 415 -3485
rect 381 -3587 415 -3553
rect 381 -3655 415 -3621
rect 381 -3723 415 -3689
rect 381 -3791 415 -3757
rect 381 -3859 415 -3825
rect 381 -3927 415 -3893
rect 381 -3995 415 -3961
rect 381 -4063 415 -4029
rect 381 -4131 415 -4097
rect 381 -4199 415 -4165
rect 381 -4267 415 -4233
rect 381 -4335 415 -4301
rect 381 -4403 415 -4369
rect 381 -4471 415 -4437
rect 381 -4539 415 -4505
rect 381 -4607 415 -4573
rect -415 -4728 -381 -4641
rect 381 -4728 415 -4641
rect -415 -4762 -289 -4728
rect -255 -4762 -221 -4728
rect -187 -4762 -153 -4728
rect -119 -4762 -85 -4728
rect -51 -4762 -17 -4728
rect 17 -4762 51 -4728
rect 85 -4762 119 -4728
rect 153 -4762 187 -4728
rect 221 -4762 255 -4728
rect 289 -4762 415 -4728
<< psubdiffcont >>
rect -289 4728 -255 4762
rect -221 4728 -187 4762
rect -153 4728 -119 4762
rect -85 4728 -51 4762
rect -17 4728 17 4762
rect 51 4728 85 4762
rect 119 4728 153 4762
rect 187 4728 221 4762
rect 255 4728 289 4762
rect -415 4607 -381 4641
rect -415 4539 -381 4573
rect -415 4471 -381 4505
rect -415 4403 -381 4437
rect -415 4335 -381 4369
rect -415 4267 -381 4301
rect -415 4199 -381 4233
rect -415 4131 -381 4165
rect -415 4063 -381 4097
rect -415 3995 -381 4029
rect -415 3927 -381 3961
rect -415 3859 -381 3893
rect -415 3791 -381 3825
rect -415 3723 -381 3757
rect -415 3655 -381 3689
rect -415 3587 -381 3621
rect -415 3519 -381 3553
rect -415 3451 -381 3485
rect -415 3383 -381 3417
rect -415 3315 -381 3349
rect -415 3247 -381 3281
rect -415 3179 -381 3213
rect -415 3111 -381 3145
rect -415 3043 -381 3077
rect -415 2975 -381 3009
rect -415 2907 -381 2941
rect -415 2839 -381 2873
rect -415 2771 -381 2805
rect -415 2703 -381 2737
rect -415 2635 -381 2669
rect -415 2567 -381 2601
rect -415 2499 -381 2533
rect -415 2431 -381 2465
rect -415 2363 -381 2397
rect -415 2295 -381 2329
rect -415 2227 -381 2261
rect -415 2159 -381 2193
rect -415 2091 -381 2125
rect -415 2023 -381 2057
rect -415 1955 -381 1989
rect -415 1887 -381 1921
rect -415 1819 -381 1853
rect -415 1751 -381 1785
rect -415 1683 -381 1717
rect -415 1615 -381 1649
rect -415 1547 -381 1581
rect -415 1479 -381 1513
rect -415 1411 -381 1445
rect -415 1343 -381 1377
rect -415 1275 -381 1309
rect -415 1207 -381 1241
rect -415 1139 -381 1173
rect -415 1071 -381 1105
rect -415 1003 -381 1037
rect -415 935 -381 969
rect -415 867 -381 901
rect -415 799 -381 833
rect -415 731 -381 765
rect -415 663 -381 697
rect -415 595 -381 629
rect -415 527 -381 561
rect -415 459 -381 493
rect -415 391 -381 425
rect -415 323 -381 357
rect -415 255 -381 289
rect -415 187 -381 221
rect -415 119 -381 153
rect -415 51 -381 85
rect -415 -17 -381 17
rect -415 -85 -381 -51
rect -415 -153 -381 -119
rect -415 -221 -381 -187
rect -415 -289 -381 -255
rect -415 -357 -381 -323
rect -415 -425 -381 -391
rect -415 -493 -381 -459
rect -415 -561 -381 -527
rect -415 -629 -381 -595
rect -415 -697 -381 -663
rect -415 -765 -381 -731
rect -415 -833 -381 -799
rect -415 -901 -381 -867
rect -415 -969 -381 -935
rect -415 -1037 -381 -1003
rect -415 -1105 -381 -1071
rect -415 -1173 -381 -1139
rect -415 -1241 -381 -1207
rect -415 -1309 -381 -1275
rect -415 -1377 -381 -1343
rect -415 -1445 -381 -1411
rect -415 -1513 -381 -1479
rect -415 -1581 -381 -1547
rect -415 -1649 -381 -1615
rect -415 -1717 -381 -1683
rect -415 -1785 -381 -1751
rect -415 -1853 -381 -1819
rect -415 -1921 -381 -1887
rect -415 -1989 -381 -1955
rect -415 -2057 -381 -2023
rect -415 -2125 -381 -2091
rect -415 -2193 -381 -2159
rect -415 -2261 -381 -2227
rect -415 -2329 -381 -2295
rect -415 -2397 -381 -2363
rect -415 -2465 -381 -2431
rect -415 -2533 -381 -2499
rect -415 -2601 -381 -2567
rect -415 -2669 -381 -2635
rect -415 -2737 -381 -2703
rect -415 -2805 -381 -2771
rect -415 -2873 -381 -2839
rect -415 -2941 -381 -2907
rect -415 -3009 -381 -2975
rect -415 -3077 -381 -3043
rect -415 -3145 -381 -3111
rect -415 -3213 -381 -3179
rect -415 -3281 -381 -3247
rect -415 -3349 -381 -3315
rect -415 -3417 -381 -3383
rect -415 -3485 -381 -3451
rect -415 -3553 -381 -3519
rect -415 -3621 -381 -3587
rect -415 -3689 -381 -3655
rect -415 -3757 -381 -3723
rect -415 -3825 -381 -3791
rect -415 -3893 -381 -3859
rect -415 -3961 -381 -3927
rect -415 -4029 -381 -3995
rect -415 -4097 -381 -4063
rect -415 -4165 -381 -4131
rect -415 -4233 -381 -4199
rect -415 -4301 -381 -4267
rect -415 -4369 -381 -4335
rect -415 -4437 -381 -4403
rect -415 -4505 -381 -4471
rect -415 -4573 -381 -4539
rect -415 -4641 -381 -4607
rect 381 4607 415 4641
rect 381 4539 415 4573
rect 381 4471 415 4505
rect 381 4403 415 4437
rect 381 4335 415 4369
rect 381 4267 415 4301
rect 381 4199 415 4233
rect 381 4131 415 4165
rect 381 4063 415 4097
rect 381 3995 415 4029
rect 381 3927 415 3961
rect 381 3859 415 3893
rect 381 3791 415 3825
rect 381 3723 415 3757
rect 381 3655 415 3689
rect 381 3587 415 3621
rect 381 3519 415 3553
rect 381 3451 415 3485
rect 381 3383 415 3417
rect 381 3315 415 3349
rect 381 3247 415 3281
rect 381 3179 415 3213
rect 381 3111 415 3145
rect 381 3043 415 3077
rect 381 2975 415 3009
rect 381 2907 415 2941
rect 381 2839 415 2873
rect 381 2771 415 2805
rect 381 2703 415 2737
rect 381 2635 415 2669
rect 381 2567 415 2601
rect 381 2499 415 2533
rect 381 2431 415 2465
rect 381 2363 415 2397
rect 381 2295 415 2329
rect 381 2227 415 2261
rect 381 2159 415 2193
rect 381 2091 415 2125
rect 381 2023 415 2057
rect 381 1955 415 1989
rect 381 1887 415 1921
rect 381 1819 415 1853
rect 381 1751 415 1785
rect 381 1683 415 1717
rect 381 1615 415 1649
rect 381 1547 415 1581
rect 381 1479 415 1513
rect 381 1411 415 1445
rect 381 1343 415 1377
rect 381 1275 415 1309
rect 381 1207 415 1241
rect 381 1139 415 1173
rect 381 1071 415 1105
rect 381 1003 415 1037
rect 381 935 415 969
rect 381 867 415 901
rect 381 799 415 833
rect 381 731 415 765
rect 381 663 415 697
rect 381 595 415 629
rect 381 527 415 561
rect 381 459 415 493
rect 381 391 415 425
rect 381 323 415 357
rect 381 255 415 289
rect 381 187 415 221
rect 381 119 415 153
rect 381 51 415 85
rect 381 -17 415 17
rect 381 -85 415 -51
rect 381 -153 415 -119
rect 381 -221 415 -187
rect 381 -289 415 -255
rect 381 -357 415 -323
rect 381 -425 415 -391
rect 381 -493 415 -459
rect 381 -561 415 -527
rect 381 -629 415 -595
rect 381 -697 415 -663
rect 381 -765 415 -731
rect 381 -833 415 -799
rect 381 -901 415 -867
rect 381 -969 415 -935
rect 381 -1037 415 -1003
rect 381 -1105 415 -1071
rect 381 -1173 415 -1139
rect 381 -1241 415 -1207
rect 381 -1309 415 -1275
rect 381 -1377 415 -1343
rect 381 -1445 415 -1411
rect 381 -1513 415 -1479
rect 381 -1581 415 -1547
rect 381 -1649 415 -1615
rect 381 -1717 415 -1683
rect 381 -1785 415 -1751
rect 381 -1853 415 -1819
rect 381 -1921 415 -1887
rect 381 -1989 415 -1955
rect 381 -2057 415 -2023
rect 381 -2125 415 -2091
rect 381 -2193 415 -2159
rect 381 -2261 415 -2227
rect 381 -2329 415 -2295
rect 381 -2397 415 -2363
rect 381 -2465 415 -2431
rect 381 -2533 415 -2499
rect 381 -2601 415 -2567
rect 381 -2669 415 -2635
rect 381 -2737 415 -2703
rect 381 -2805 415 -2771
rect 381 -2873 415 -2839
rect 381 -2941 415 -2907
rect 381 -3009 415 -2975
rect 381 -3077 415 -3043
rect 381 -3145 415 -3111
rect 381 -3213 415 -3179
rect 381 -3281 415 -3247
rect 381 -3349 415 -3315
rect 381 -3417 415 -3383
rect 381 -3485 415 -3451
rect 381 -3553 415 -3519
rect 381 -3621 415 -3587
rect 381 -3689 415 -3655
rect 381 -3757 415 -3723
rect 381 -3825 415 -3791
rect 381 -3893 415 -3859
rect 381 -3961 415 -3927
rect 381 -4029 415 -3995
rect 381 -4097 415 -4063
rect 381 -4165 415 -4131
rect 381 -4233 415 -4199
rect 381 -4301 415 -4267
rect 381 -4369 415 -4335
rect 381 -4437 415 -4403
rect 381 -4505 415 -4471
rect 381 -4573 415 -4539
rect 381 -4641 415 -4607
rect -289 -4762 -255 -4728
rect -221 -4762 -187 -4728
rect -153 -4762 -119 -4728
rect -85 -4762 -51 -4728
rect -17 -4762 17 -4728
rect 51 -4762 85 -4728
rect 119 -4762 153 -4728
rect 187 -4762 221 -4728
rect 255 -4762 289 -4728
<< xpolycontact >>
rect -285 4200 285 4632
rect -285 -4632 285 -4200
<< ppolyres >>
rect -285 -4200 285 4200
<< locali >>
rect -415 4728 -289 4762
rect -255 4728 -221 4762
rect -187 4728 -153 4762
rect -119 4728 -85 4762
rect -51 4728 -17 4762
rect 17 4728 51 4762
rect 85 4728 119 4762
rect 153 4728 187 4762
rect 221 4728 255 4762
rect 289 4728 415 4762
rect -415 4641 -381 4728
rect 381 4641 415 4728
rect -415 4573 -381 4607
rect -415 4505 -381 4539
rect -415 4437 -381 4471
rect -415 4369 -381 4403
rect -415 4301 -381 4335
rect -415 4233 -381 4267
rect 381 4573 415 4607
rect 381 4505 415 4539
rect 381 4437 415 4471
rect 381 4369 415 4403
rect 381 4301 415 4335
rect 381 4233 415 4267
rect -415 4165 -381 4199
rect -415 4097 -381 4131
rect -415 4029 -381 4063
rect -415 3961 -381 3995
rect -415 3893 -381 3927
rect -415 3825 -381 3859
rect -415 3757 -381 3791
rect -415 3689 -381 3723
rect -415 3621 -381 3655
rect -415 3553 -381 3587
rect -415 3485 -381 3519
rect -415 3417 -381 3451
rect -415 3349 -381 3383
rect -415 3281 -381 3315
rect -415 3213 -381 3247
rect -415 3145 -381 3179
rect -415 3077 -381 3111
rect -415 3009 -381 3043
rect -415 2941 -381 2975
rect -415 2873 -381 2907
rect -415 2805 -381 2839
rect -415 2737 -381 2771
rect -415 2669 -381 2703
rect -415 2601 -381 2635
rect -415 2533 -381 2567
rect -415 2465 -381 2499
rect -415 2397 -381 2431
rect -415 2329 -381 2363
rect -415 2261 -381 2295
rect -415 2193 -381 2227
rect -415 2125 -381 2159
rect -415 2057 -381 2091
rect -415 1989 -381 2023
rect -415 1921 -381 1955
rect -415 1853 -381 1887
rect -415 1785 -381 1819
rect -415 1717 -381 1751
rect -415 1649 -381 1683
rect -415 1581 -381 1615
rect -415 1513 -381 1547
rect -415 1445 -381 1479
rect -415 1377 -381 1411
rect -415 1309 -381 1343
rect -415 1241 -381 1275
rect -415 1173 -381 1207
rect -415 1105 -381 1139
rect -415 1037 -381 1071
rect -415 969 -381 1003
rect -415 901 -381 935
rect -415 833 -381 867
rect -415 765 -381 799
rect -415 697 -381 731
rect -415 629 -381 663
rect -415 561 -381 595
rect -415 493 -381 527
rect -415 425 -381 459
rect -415 357 -381 391
rect -415 289 -381 323
rect -415 221 -381 255
rect -415 153 -381 187
rect -415 85 -381 119
rect -415 17 -381 51
rect -415 -51 -381 -17
rect -415 -119 -381 -85
rect -415 -187 -381 -153
rect -415 -255 -381 -221
rect -415 -323 -381 -289
rect -415 -391 -381 -357
rect -415 -459 -381 -425
rect -415 -527 -381 -493
rect -415 -595 -381 -561
rect -415 -663 -381 -629
rect -415 -731 -381 -697
rect -415 -799 -381 -765
rect -415 -867 -381 -833
rect -415 -935 -381 -901
rect -415 -1003 -381 -969
rect -415 -1071 -381 -1037
rect -415 -1139 -381 -1105
rect -415 -1207 -381 -1173
rect -415 -1275 -381 -1241
rect -415 -1343 -381 -1309
rect -415 -1411 -381 -1377
rect -415 -1479 -381 -1445
rect -415 -1547 -381 -1513
rect -415 -1615 -381 -1581
rect -415 -1683 -381 -1649
rect -415 -1751 -381 -1717
rect -415 -1819 -381 -1785
rect -415 -1887 -381 -1853
rect -415 -1955 -381 -1921
rect -415 -2023 -381 -1989
rect -415 -2091 -381 -2057
rect -415 -2159 -381 -2125
rect -415 -2227 -381 -2193
rect -415 -2295 -381 -2261
rect -415 -2363 -381 -2329
rect -415 -2431 -381 -2397
rect -415 -2499 -381 -2465
rect -415 -2567 -381 -2533
rect -415 -2635 -381 -2601
rect -415 -2703 -381 -2669
rect -415 -2771 -381 -2737
rect -415 -2839 -381 -2805
rect -415 -2907 -381 -2873
rect -415 -2975 -381 -2941
rect -415 -3043 -381 -3009
rect -415 -3111 -381 -3077
rect -415 -3179 -381 -3145
rect -415 -3247 -381 -3213
rect -415 -3315 -381 -3281
rect -415 -3383 -381 -3349
rect -415 -3451 -381 -3417
rect -415 -3519 -381 -3485
rect -415 -3587 -381 -3553
rect -415 -3655 -381 -3621
rect -415 -3723 -381 -3689
rect -415 -3791 -381 -3757
rect -415 -3859 -381 -3825
rect -415 -3927 -381 -3893
rect -415 -3995 -381 -3961
rect -415 -4063 -381 -4029
rect -415 -4131 -381 -4097
rect -415 -4199 -381 -4165
rect 381 4165 415 4199
rect 381 4097 415 4131
rect 381 4029 415 4063
rect 381 3961 415 3995
rect 381 3893 415 3927
rect 381 3825 415 3859
rect 381 3757 415 3791
rect 381 3689 415 3723
rect 381 3621 415 3655
rect 381 3553 415 3587
rect 381 3485 415 3519
rect 381 3417 415 3451
rect 381 3349 415 3383
rect 381 3281 415 3315
rect 381 3213 415 3247
rect 381 3145 415 3179
rect 381 3077 415 3111
rect 381 3009 415 3043
rect 381 2941 415 2975
rect 381 2873 415 2907
rect 381 2805 415 2839
rect 381 2737 415 2771
rect 381 2669 415 2703
rect 381 2601 415 2635
rect 381 2533 415 2567
rect 381 2465 415 2499
rect 381 2397 415 2431
rect 381 2329 415 2363
rect 381 2261 415 2295
rect 381 2193 415 2227
rect 381 2125 415 2159
rect 381 2057 415 2091
rect 381 1989 415 2023
rect 381 1921 415 1955
rect 381 1853 415 1887
rect 381 1785 415 1819
rect 381 1717 415 1751
rect 381 1649 415 1683
rect 381 1581 415 1615
rect 381 1513 415 1547
rect 381 1445 415 1479
rect 381 1377 415 1411
rect 381 1309 415 1343
rect 381 1241 415 1275
rect 381 1173 415 1207
rect 381 1105 415 1139
rect 381 1037 415 1071
rect 381 969 415 1003
rect 381 901 415 935
rect 381 833 415 867
rect 381 765 415 799
rect 381 697 415 731
rect 381 629 415 663
rect 381 561 415 595
rect 381 493 415 527
rect 381 425 415 459
rect 381 357 415 391
rect 381 289 415 323
rect 381 221 415 255
rect 381 153 415 187
rect 381 85 415 119
rect 381 17 415 51
rect 381 -51 415 -17
rect 381 -119 415 -85
rect 381 -187 415 -153
rect 381 -255 415 -221
rect 381 -323 415 -289
rect 381 -391 415 -357
rect 381 -459 415 -425
rect 381 -527 415 -493
rect 381 -595 415 -561
rect 381 -663 415 -629
rect 381 -731 415 -697
rect 381 -799 415 -765
rect 381 -867 415 -833
rect 381 -935 415 -901
rect 381 -1003 415 -969
rect 381 -1071 415 -1037
rect 381 -1139 415 -1105
rect 381 -1207 415 -1173
rect 381 -1275 415 -1241
rect 381 -1343 415 -1309
rect 381 -1411 415 -1377
rect 381 -1479 415 -1445
rect 381 -1547 415 -1513
rect 381 -1615 415 -1581
rect 381 -1683 415 -1649
rect 381 -1751 415 -1717
rect 381 -1819 415 -1785
rect 381 -1887 415 -1853
rect 381 -1955 415 -1921
rect 381 -2023 415 -1989
rect 381 -2091 415 -2057
rect 381 -2159 415 -2125
rect 381 -2227 415 -2193
rect 381 -2295 415 -2261
rect 381 -2363 415 -2329
rect 381 -2431 415 -2397
rect 381 -2499 415 -2465
rect 381 -2567 415 -2533
rect 381 -2635 415 -2601
rect 381 -2703 415 -2669
rect 381 -2771 415 -2737
rect 381 -2839 415 -2805
rect 381 -2907 415 -2873
rect 381 -2975 415 -2941
rect 381 -3043 415 -3009
rect 381 -3111 415 -3077
rect 381 -3179 415 -3145
rect 381 -3247 415 -3213
rect 381 -3315 415 -3281
rect 381 -3383 415 -3349
rect 381 -3451 415 -3417
rect 381 -3519 415 -3485
rect 381 -3587 415 -3553
rect 381 -3655 415 -3621
rect 381 -3723 415 -3689
rect 381 -3791 415 -3757
rect 381 -3859 415 -3825
rect 381 -3927 415 -3893
rect 381 -3995 415 -3961
rect 381 -4063 415 -4029
rect 381 -4131 415 -4097
rect 381 -4199 415 -4165
rect -415 -4267 -381 -4233
rect -415 -4335 -381 -4301
rect -415 -4403 -381 -4369
rect -415 -4471 -381 -4437
rect -415 -4539 -381 -4505
rect -415 -4607 -381 -4573
rect 381 -4267 415 -4233
rect 381 -4335 415 -4301
rect 381 -4403 415 -4369
rect 381 -4471 415 -4437
rect 381 -4539 415 -4505
rect 381 -4607 415 -4573
rect -415 -4728 -381 -4641
rect 381 -4728 415 -4641
rect -415 -4762 -289 -4728
rect -255 -4762 -221 -4728
rect -187 -4762 -153 -4728
rect -119 -4762 -85 -4728
rect -51 -4762 -17 -4728
rect 17 -4762 51 -4728
rect 85 -4762 119 -4728
rect 153 -4762 187 -4728
rect 221 -4762 255 -4728
rect 289 -4762 415 -4728
<< viali >>
rect -269 4218 269 4612
rect -269 -4613 269 -4219
<< metal1 >>
rect -281 4612 281 4620
rect -281 4218 -269 4612
rect 269 4218 281 4612
rect -281 4211 281 4218
rect -281 -4219 281 -4211
rect -281 -4613 -269 -4219
rect 269 -4613 281 -4219
rect -281 -4620 281 -4613
<< properties >>
string FIXED_BBOX -398 -4745 398 4745
<< end >>
