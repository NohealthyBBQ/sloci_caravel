magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect -17320 14867 35240 14880
rect -17320 14833 -17301 14867
rect -17267 14833 -17229 14867
rect -17195 14833 -17157 14867
rect -17123 14833 -17085 14867
rect -17051 14833 -17013 14867
rect -16979 14833 -16941 14867
rect -16907 14833 -16869 14867
rect -16835 14833 -16797 14867
rect -16763 14833 -16725 14867
rect -16691 14833 -16653 14867
rect -16619 14833 -16581 14867
rect -16547 14833 -16509 14867
rect -16475 14833 -16437 14867
rect -16403 14833 -16365 14867
rect -16331 14833 -16293 14867
rect -16259 14833 -16221 14867
rect -16187 14833 -16149 14867
rect -16115 14833 -16077 14867
rect -16043 14833 -16005 14867
rect -15971 14833 -15933 14867
rect -15899 14833 -15861 14867
rect -15827 14833 -15789 14867
rect -15755 14833 -15717 14867
rect -15683 14833 -15645 14867
rect -15611 14833 -15573 14867
rect -15539 14833 -15501 14867
rect -15467 14833 -15429 14867
rect -15395 14833 -15357 14867
rect -15323 14833 -15285 14867
rect -15251 14833 -15213 14867
rect -15179 14833 -15141 14867
rect -15107 14833 -15069 14867
rect -15035 14833 -14997 14867
rect -14963 14833 -14925 14867
rect -14891 14833 -14853 14867
rect -14819 14833 -14781 14867
rect -14747 14833 -14709 14867
rect -14675 14833 -14637 14867
rect -14603 14833 -14565 14867
rect -14531 14833 -14493 14867
rect -14459 14833 -14421 14867
rect -14387 14833 -14349 14867
rect -14315 14833 -14277 14867
rect -14243 14833 -14205 14867
rect -14171 14833 -14133 14867
rect -14099 14833 -14061 14867
rect -14027 14833 -13989 14867
rect -13955 14833 -13917 14867
rect -13883 14833 -13845 14867
rect -13811 14833 -13773 14867
rect -13739 14833 -13701 14867
rect -13667 14833 -13629 14867
rect -13595 14833 -13557 14867
rect -13523 14833 -13485 14867
rect -13451 14833 -13413 14867
rect -13379 14833 -13341 14867
rect -13307 14833 -13269 14867
rect -13235 14833 -13197 14867
rect -13163 14833 -13125 14867
rect -13091 14833 -13053 14867
rect -13019 14833 -12981 14867
rect -12947 14833 -12909 14867
rect -12875 14833 -12837 14867
rect -12803 14833 -12765 14867
rect -12731 14833 -12693 14867
rect -12659 14833 -12621 14867
rect -12587 14833 -12549 14867
rect -12515 14833 -12477 14867
rect -12443 14833 -12405 14867
rect -12371 14833 -12333 14867
rect -12299 14833 -12261 14867
rect -12227 14833 -12189 14867
rect -12155 14833 -12117 14867
rect -12083 14833 -12045 14867
rect -12011 14833 -11973 14867
rect -11939 14833 -11901 14867
rect -11867 14833 -11829 14867
rect -11795 14833 -11757 14867
rect -11723 14833 -11685 14867
rect -11651 14833 -11613 14867
rect -11579 14833 -11541 14867
rect -11507 14833 -11469 14867
rect -11435 14833 -11397 14867
rect -11363 14833 -11325 14867
rect -11291 14833 -11253 14867
rect -11219 14833 -11181 14867
rect -11147 14833 -11109 14867
rect -11075 14833 -11037 14867
rect -11003 14833 -10965 14867
rect -10931 14833 -10893 14867
rect -10859 14833 -10821 14867
rect -10787 14833 -10749 14867
rect -10715 14833 -10677 14867
rect -10643 14833 -10605 14867
rect -10571 14833 -10533 14867
rect -10499 14833 -10461 14867
rect -10427 14833 -10389 14867
rect -10355 14833 -10317 14867
rect -10283 14833 -10245 14867
rect -10211 14833 -10173 14867
rect -10139 14833 -10101 14867
rect -10067 14833 -10029 14867
rect -9995 14833 -9957 14867
rect -9923 14833 -9885 14867
rect -9851 14833 -9813 14867
rect -9779 14833 -9741 14867
rect -9707 14833 -9669 14867
rect -9635 14833 -9597 14867
rect -9563 14833 -9525 14867
rect -9491 14833 -9453 14867
rect -9419 14833 -9381 14867
rect -9347 14833 -9309 14867
rect -9275 14833 -9237 14867
rect -9203 14833 -9165 14867
rect -9131 14833 -9093 14867
rect -9059 14833 -9021 14867
rect -8987 14833 -8949 14867
rect -8915 14833 -8877 14867
rect -8843 14833 -8805 14867
rect -8771 14833 -8733 14867
rect -8699 14833 -8661 14867
rect -8627 14833 -8589 14867
rect -8555 14833 -8517 14867
rect -8483 14833 -8445 14867
rect -8411 14833 -8373 14867
rect -8339 14833 -8301 14867
rect -8267 14833 -8229 14867
rect -8195 14833 -8157 14867
rect -8123 14833 -8085 14867
rect -8051 14833 -8013 14867
rect -7979 14833 -7941 14867
rect -7907 14833 -7869 14867
rect -7835 14833 -7797 14867
rect -7763 14833 -7725 14867
rect -7691 14833 -7653 14867
rect -7619 14833 -7581 14867
rect -7547 14833 -7509 14867
rect -7475 14833 -7437 14867
rect -7403 14833 -7365 14867
rect -7331 14833 -7293 14867
rect -7259 14833 -7221 14867
rect -7187 14833 -7149 14867
rect -7115 14833 -7077 14867
rect -7043 14833 -7005 14867
rect -6971 14833 -6933 14867
rect -6899 14833 -6861 14867
rect -6827 14833 -6789 14867
rect -6755 14833 -6717 14867
rect -6683 14833 -6645 14867
rect -6611 14833 -6573 14867
rect -6539 14833 -6501 14867
rect -6467 14833 -6429 14867
rect -6395 14833 -6357 14867
rect -6323 14833 -6285 14867
rect -6251 14833 -6213 14867
rect -6179 14833 -6141 14867
rect -6107 14833 -6069 14867
rect -6035 14833 -5997 14867
rect -5963 14833 -5925 14867
rect -5891 14833 -5853 14867
rect -5819 14833 -5781 14867
rect -5747 14833 -5709 14867
rect -5675 14833 -5637 14867
rect -5603 14833 -5565 14867
rect -5531 14833 -5493 14867
rect -5459 14833 -5421 14867
rect -5387 14833 -5349 14867
rect -5315 14833 -5277 14867
rect -5243 14833 -5205 14867
rect -5171 14833 -5133 14867
rect -5099 14833 -5061 14867
rect -5027 14833 -4989 14867
rect -4955 14833 -4917 14867
rect -4883 14833 -4845 14867
rect -4811 14833 -4773 14867
rect -4739 14833 -4701 14867
rect -4667 14833 -4629 14867
rect -4595 14833 -4557 14867
rect -4523 14833 -4485 14867
rect -4451 14833 -4413 14867
rect -4379 14833 -4341 14867
rect -4307 14833 -4269 14867
rect -4235 14833 -4197 14867
rect -4163 14833 -4125 14867
rect -4091 14833 -4053 14867
rect -4019 14833 -3981 14867
rect -3947 14833 -3909 14867
rect -3875 14833 -3837 14867
rect -3803 14833 -3765 14867
rect -3731 14833 -3693 14867
rect -3659 14833 -3621 14867
rect -3587 14833 -3549 14867
rect -3515 14833 -3477 14867
rect -3443 14833 -3405 14867
rect -3371 14833 -3333 14867
rect -3299 14833 -3261 14867
rect -3227 14833 -3189 14867
rect -3155 14833 -3117 14867
rect -3083 14833 -3045 14867
rect -3011 14833 -2973 14867
rect -2939 14833 -2901 14867
rect -2867 14833 -2829 14867
rect -2795 14833 -2757 14867
rect -2723 14833 -2685 14867
rect -2651 14833 -2613 14867
rect -2579 14833 -2541 14867
rect -2507 14833 -2469 14867
rect -2435 14833 -2397 14867
rect -2363 14833 -2325 14867
rect -2291 14833 -2253 14867
rect -2219 14833 -2181 14867
rect -2147 14833 -2109 14867
rect -2075 14833 -2037 14867
rect -2003 14833 -1965 14867
rect -1931 14833 -1893 14867
rect -1859 14833 -1821 14867
rect -1787 14833 -1749 14867
rect -1715 14833 -1677 14867
rect -1643 14833 -1605 14867
rect -1571 14833 -1533 14867
rect -1499 14833 -1461 14867
rect -1427 14833 -1389 14867
rect -1355 14833 -1317 14867
rect -1283 14833 -1245 14867
rect -1211 14833 -1173 14867
rect -1139 14833 -1101 14867
rect -1067 14833 -1029 14867
rect -995 14833 -957 14867
rect -923 14833 -885 14867
rect -851 14833 -813 14867
rect -779 14833 -741 14867
rect -707 14833 -669 14867
rect -635 14833 -597 14867
rect -563 14833 -525 14867
rect -491 14833 -453 14867
rect -419 14833 -381 14867
rect -347 14833 -309 14867
rect -275 14833 -237 14867
rect -203 14833 -165 14867
rect -131 14833 -93 14867
rect -59 14833 -21 14867
rect 13 14833 51 14867
rect 85 14833 123 14867
rect 157 14833 195 14867
rect 229 14833 267 14867
rect 301 14833 339 14867
rect 373 14833 411 14867
rect 445 14833 483 14867
rect 517 14833 555 14867
rect 589 14833 627 14867
rect 661 14833 699 14867
rect 733 14833 771 14867
rect 805 14833 843 14867
rect 877 14833 915 14867
rect 949 14833 987 14867
rect 1021 14833 1059 14867
rect 1093 14833 1131 14867
rect 1165 14833 1203 14867
rect 1237 14833 1275 14867
rect 1309 14833 1347 14867
rect 1381 14833 1419 14867
rect 1453 14833 1491 14867
rect 1525 14833 1563 14867
rect 1597 14833 1635 14867
rect 1669 14833 1707 14867
rect 1741 14833 1779 14867
rect 1813 14833 1851 14867
rect 1885 14833 1923 14867
rect 1957 14833 1995 14867
rect 2029 14833 2067 14867
rect 2101 14833 2139 14867
rect 2173 14833 2211 14867
rect 2245 14833 2283 14867
rect 2317 14833 2355 14867
rect 2389 14833 2427 14867
rect 2461 14833 2499 14867
rect 2533 14833 2571 14867
rect 2605 14833 2643 14867
rect 2677 14833 2715 14867
rect 2749 14833 2787 14867
rect 2821 14833 2859 14867
rect 2893 14833 2931 14867
rect 2965 14833 3003 14867
rect 3037 14833 3075 14867
rect 3109 14833 3147 14867
rect 3181 14833 3219 14867
rect 3253 14833 3291 14867
rect 3325 14833 3363 14867
rect 3397 14833 3435 14867
rect 3469 14833 3507 14867
rect 3541 14833 3579 14867
rect 3613 14833 3651 14867
rect 3685 14833 3723 14867
rect 3757 14833 3795 14867
rect 3829 14833 3867 14867
rect 3901 14833 3939 14867
rect 3973 14833 4011 14867
rect 4045 14833 4083 14867
rect 4117 14833 4155 14867
rect 4189 14833 4227 14867
rect 4261 14833 4299 14867
rect 4333 14833 4371 14867
rect 4405 14833 4443 14867
rect 4477 14833 4515 14867
rect 4549 14833 4587 14867
rect 4621 14833 4659 14867
rect 4693 14833 4731 14867
rect 4765 14833 4803 14867
rect 4837 14833 4875 14867
rect 4909 14833 4947 14867
rect 4981 14833 5019 14867
rect 5053 14833 5091 14867
rect 5125 14833 5163 14867
rect 5197 14833 5235 14867
rect 5269 14833 5307 14867
rect 5341 14833 5379 14867
rect 5413 14833 5451 14867
rect 5485 14833 5523 14867
rect 5557 14833 5595 14867
rect 5629 14833 5667 14867
rect 5701 14833 5739 14867
rect 5773 14833 5811 14867
rect 5845 14833 5883 14867
rect 5917 14833 5955 14867
rect 5989 14833 6027 14867
rect 6061 14833 6099 14867
rect 6133 14833 6171 14867
rect 6205 14833 6243 14867
rect 6277 14833 6315 14867
rect 6349 14833 6387 14867
rect 6421 14833 6459 14867
rect 6493 14833 6531 14867
rect 6565 14833 6603 14867
rect 6637 14833 6675 14867
rect 6709 14833 6747 14867
rect 6781 14833 6819 14867
rect 6853 14833 6891 14867
rect 6925 14833 6963 14867
rect 6997 14833 7035 14867
rect 7069 14833 7107 14867
rect 7141 14833 7179 14867
rect 7213 14833 7251 14867
rect 7285 14833 7323 14867
rect 7357 14833 7395 14867
rect 7429 14833 7467 14867
rect 7501 14833 7539 14867
rect 7573 14833 7611 14867
rect 7645 14833 7683 14867
rect 7717 14833 7755 14867
rect 7789 14833 7827 14867
rect 7861 14833 7899 14867
rect 7933 14833 7971 14867
rect 8005 14833 8043 14867
rect 8077 14833 8115 14867
rect 8149 14833 8187 14867
rect 8221 14833 8259 14867
rect 8293 14833 8331 14867
rect 8365 14833 8403 14867
rect 8437 14833 8475 14867
rect 8509 14833 8547 14867
rect 8581 14833 8619 14867
rect 8653 14833 8691 14867
rect 8725 14833 8763 14867
rect 8797 14833 8835 14867
rect 8869 14833 8907 14867
rect 8941 14833 8979 14867
rect 9013 14833 9051 14867
rect 9085 14833 9123 14867
rect 9157 14833 9195 14867
rect 9229 14833 9267 14867
rect 9301 14833 9339 14867
rect 9373 14833 9411 14867
rect 9445 14833 9483 14867
rect 9517 14833 9555 14867
rect 9589 14833 9627 14867
rect 9661 14833 9699 14867
rect 9733 14833 9771 14867
rect 9805 14833 9843 14867
rect 9877 14833 9915 14867
rect 9949 14833 9987 14867
rect 10021 14833 10059 14867
rect 10093 14833 10131 14867
rect 10165 14833 10203 14867
rect 10237 14833 10275 14867
rect 10309 14833 10347 14867
rect 10381 14833 10419 14867
rect 10453 14833 10491 14867
rect 10525 14833 10563 14867
rect 10597 14833 10635 14867
rect 10669 14833 10707 14867
rect 10741 14833 10779 14867
rect 10813 14833 10851 14867
rect 10885 14833 10923 14867
rect 10957 14833 10995 14867
rect 11029 14833 11067 14867
rect 11101 14833 11139 14867
rect 11173 14833 11211 14867
rect 11245 14833 11283 14867
rect 11317 14833 11355 14867
rect 11389 14833 11427 14867
rect 11461 14833 11499 14867
rect 11533 14833 11571 14867
rect 11605 14833 11643 14867
rect 11677 14833 11715 14867
rect 11749 14833 11787 14867
rect 11821 14833 11859 14867
rect 11893 14833 11931 14867
rect 11965 14833 12003 14867
rect 12037 14833 12075 14867
rect 12109 14833 12147 14867
rect 12181 14833 12219 14867
rect 12253 14833 12291 14867
rect 12325 14833 12363 14867
rect 12397 14833 12435 14867
rect 12469 14833 12507 14867
rect 12541 14833 12579 14867
rect 12613 14833 12651 14867
rect 12685 14833 12723 14867
rect 12757 14833 12795 14867
rect 12829 14833 12867 14867
rect 12901 14833 12939 14867
rect 12973 14833 13011 14867
rect 13045 14833 13083 14867
rect 13117 14833 13155 14867
rect 13189 14833 13227 14867
rect 13261 14833 13299 14867
rect 13333 14833 13371 14867
rect 13405 14833 13443 14867
rect 13477 14833 13515 14867
rect 13549 14833 13587 14867
rect 13621 14833 13659 14867
rect 13693 14833 13731 14867
rect 13765 14833 13803 14867
rect 13837 14833 13875 14867
rect 13909 14833 13947 14867
rect 13981 14833 14019 14867
rect 14053 14833 14091 14867
rect 14125 14833 14163 14867
rect 14197 14833 14235 14867
rect 14269 14833 14307 14867
rect 14341 14833 14379 14867
rect 14413 14833 14451 14867
rect 14485 14833 14523 14867
rect 14557 14833 14595 14867
rect 14629 14833 14667 14867
rect 14701 14833 14739 14867
rect 14773 14833 14811 14867
rect 14845 14833 14883 14867
rect 14917 14833 14955 14867
rect 14989 14833 15027 14867
rect 15061 14833 15099 14867
rect 15133 14833 15171 14867
rect 15205 14833 15243 14867
rect 15277 14833 15315 14867
rect 15349 14833 15387 14867
rect 15421 14833 15459 14867
rect 15493 14833 15531 14867
rect 15565 14833 15603 14867
rect 15637 14833 15675 14867
rect 15709 14833 15747 14867
rect 15781 14833 15819 14867
rect 15853 14833 15891 14867
rect 15925 14833 15963 14867
rect 15997 14833 16035 14867
rect 16069 14833 16107 14867
rect 16141 14833 16179 14867
rect 16213 14833 16251 14867
rect 16285 14833 16323 14867
rect 16357 14833 16395 14867
rect 16429 14833 16467 14867
rect 16501 14833 16539 14867
rect 16573 14833 16611 14867
rect 16645 14833 16683 14867
rect 16717 14833 16755 14867
rect 16789 14833 16827 14867
rect 16861 14833 16899 14867
rect 16933 14833 16971 14867
rect 17005 14833 17043 14867
rect 17077 14833 17115 14867
rect 17149 14833 17187 14867
rect 17221 14833 17259 14867
rect 17293 14833 17331 14867
rect 17365 14833 17403 14867
rect 17437 14833 17475 14867
rect 17509 14833 17547 14867
rect 17581 14833 17619 14867
rect 17653 14833 17691 14867
rect 17725 14833 17763 14867
rect 17797 14833 17835 14867
rect 17869 14833 17907 14867
rect 17941 14833 17979 14867
rect 18013 14833 18051 14867
rect 18085 14833 18123 14867
rect 18157 14833 18195 14867
rect 18229 14833 18267 14867
rect 18301 14833 18339 14867
rect 18373 14833 18411 14867
rect 18445 14833 18483 14867
rect 18517 14833 18555 14867
rect 18589 14833 18627 14867
rect 18661 14833 18699 14867
rect 18733 14833 18771 14867
rect 18805 14833 18843 14867
rect 18877 14833 18915 14867
rect 18949 14833 18987 14867
rect 19021 14833 19059 14867
rect 19093 14833 19131 14867
rect 19165 14833 19203 14867
rect 19237 14833 19275 14867
rect 19309 14833 19347 14867
rect 19381 14833 19419 14867
rect 19453 14833 19491 14867
rect 19525 14833 19563 14867
rect 19597 14833 19635 14867
rect 19669 14833 19707 14867
rect 19741 14833 19779 14867
rect 19813 14833 19851 14867
rect 19885 14833 19923 14867
rect 19957 14833 19995 14867
rect 20029 14833 20067 14867
rect 20101 14833 20139 14867
rect 20173 14833 20211 14867
rect 20245 14833 20283 14867
rect 20317 14833 20355 14867
rect 20389 14833 20427 14867
rect 20461 14833 20499 14867
rect 20533 14833 20571 14867
rect 20605 14833 20643 14867
rect 20677 14833 20715 14867
rect 20749 14833 20787 14867
rect 20821 14833 20859 14867
rect 20893 14833 20931 14867
rect 20965 14833 21003 14867
rect 21037 14833 21075 14867
rect 21109 14833 21147 14867
rect 21181 14833 21219 14867
rect 21253 14833 21291 14867
rect 21325 14833 21363 14867
rect 21397 14833 21435 14867
rect 21469 14833 21507 14867
rect 21541 14833 21579 14867
rect 21613 14833 21651 14867
rect 21685 14833 21723 14867
rect 21757 14833 21795 14867
rect 21829 14833 21867 14867
rect 21901 14833 21939 14867
rect 21973 14833 22011 14867
rect 22045 14833 22083 14867
rect 22117 14833 22155 14867
rect 22189 14833 22227 14867
rect 22261 14833 22299 14867
rect 22333 14833 22371 14867
rect 22405 14833 22443 14867
rect 22477 14833 22515 14867
rect 22549 14833 22587 14867
rect 22621 14833 22659 14867
rect 22693 14833 22731 14867
rect 22765 14833 22803 14867
rect 22837 14833 22875 14867
rect 22909 14833 22947 14867
rect 22981 14833 23019 14867
rect 23053 14833 23091 14867
rect 23125 14833 23163 14867
rect 23197 14833 23235 14867
rect 23269 14833 23307 14867
rect 23341 14833 23379 14867
rect 23413 14833 23451 14867
rect 23485 14833 23523 14867
rect 23557 14833 23595 14867
rect 23629 14833 23667 14867
rect 23701 14833 23739 14867
rect 23773 14833 23811 14867
rect 23845 14833 23883 14867
rect 23917 14833 23955 14867
rect 23989 14833 24027 14867
rect 24061 14833 24099 14867
rect 24133 14833 24171 14867
rect 24205 14833 24243 14867
rect 24277 14833 24315 14867
rect 24349 14833 24387 14867
rect 24421 14833 24459 14867
rect 24493 14833 24531 14867
rect 24565 14833 24603 14867
rect 24637 14833 24675 14867
rect 24709 14833 24747 14867
rect 24781 14833 24819 14867
rect 24853 14833 24891 14867
rect 24925 14833 24963 14867
rect 24997 14833 25035 14867
rect 25069 14833 25107 14867
rect 25141 14833 25179 14867
rect 25213 14833 25251 14867
rect 25285 14833 25323 14867
rect 25357 14833 25395 14867
rect 25429 14833 25467 14867
rect 25501 14833 25539 14867
rect 25573 14833 25611 14867
rect 25645 14833 25683 14867
rect 25717 14833 25755 14867
rect 25789 14833 25827 14867
rect 25861 14833 25899 14867
rect 25933 14833 25971 14867
rect 26005 14833 26043 14867
rect 26077 14833 26115 14867
rect 26149 14833 26187 14867
rect 26221 14833 26259 14867
rect 26293 14833 26331 14867
rect 26365 14833 26403 14867
rect 26437 14833 26475 14867
rect 26509 14833 26547 14867
rect 26581 14833 26619 14867
rect 26653 14833 26691 14867
rect 26725 14833 26763 14867
rect 26797 14833 26835 14867
rect 26869 14833 26907 14867
rect 26941 14833 26979 14867
rect 27013 14833 27051 14867
rect 27085 14833 27123 14867
rect 27157 14833 27195 14867
rect 27229 14833 27267 14867
rect 27301 14833 27339 14867
rect 27373 14833 27411 14867
rect 27445 14833 27483 14867
rect 27517 14833 27555 14867
rect 27589 14833 27627 14867
rect 27661 14833 27699 14867
rect 27733 14833 27771 14867
rect 27805 14833 27843 14867
rect 27877 14833 27915 14867
rect 27949 14833 27987 14867
rect 28021 14833 28059 14867
rect 28093 14833 28131 14867
rect 28165 14833 28203 14867
rect 28237 14833 28275 14867
rect 28309 14833 28347 14867
rect 28381 14833 28419 14867
rect 28453 14833 28491 14867
rect 28525 14833 28563 14867
rect 28597 14833 28635 14867
rect 28669 14833 28707 14867
rect 28741 14833 28779 14867
rect 28813 14833 28851 14867
rect 28885 14833 28923 14867
rect 28957 14833 28995 14867
rect 29029 14833 29067 14867
rect 29101 14833 29139 14867
rect 29173 14833 29211 14867
rect 29245 14833 29283 14867
rect 29317 14833 29355 14867
rect 29389 14833 29427 14867
rect 29461 14833 29499 14867
rect 29533 14833 29571 14867
rect 29605 14833 29643 14867
rect 29677 14833 29715 14867
rect 29749 14833 29787 14867
rect 29821 14833 29859 14867
rect 29893 14833 29931 14867
rect 29965 14833 30003 14867
rect 30037 14833 30075 14867
rect 30109 14833 30147 14867
rect 30181 14833 30219 14867
rect 30253 14833 30291 14867
rect 30325 14833 30363 14867
rect 30397 14833 30435 14867
rect 30469 14833 30507 14867
rect 30541 14833 30579 14867
rect 30613 14833 30651 14867
rect 30685 14833 30723 14867
rect 30757 14833 30795 14867
rect 30829 14833 30867 14867
rect 30901 14833 30939 14867
rect 30973 14833 31011 14867
rect 31045 14833 31083 14867
rect 31117 14833 31155 14867
rect 31189 14833 31227 14867
rect 31261 14833 31299 14867
rect 31333 14833 31371 14867
rect 31405 14833 31443 14867
rect 31477 14833 31515 14867
rect 31549 14833 31587 14867
rect 31621 14833 31659 14867
rect 31693 14833 31731 14867
rect 31765 14833 31803 14867
rect 31837 14833 31875 14867
rect 31909 14833 31947 14867
rect 31981 14833 32019 14867
rect 32053 14833 32091 14867
rect 32125 14833 32163 14867
rect 32197 14833 32235 14867
rect 32269 14833 32307 14867
rect 32341 14833 32379 14867
rect 32413 14833 32451 14867
rect 32485 14833 32523 14867
rect 32557 14833 32595 14867
rect 32629 14833 32667 14867
rect 32701 14833 32739 14867
rect 32773 14833 32811 14867
rect 32845 14833 32883 14867
rect 32917 14833 32955 14867
rect 32989 14833 33027 14867
rect 33061 14833 33099 14867
rect 33133 14833 33171 14867
rect 33205 14833 33243 14867
rect 33277 14833 33315 14867
rect 33349 14833 33387 14867
rect 33421 14833 33459 14867
rect 33493 14833 33531 14867
rect 33565 14833 33603 14867
rect 33637 14833 33675 14867
rect 33709 14833 33747 14867
rect 33781 14833 33819 14867
rect 33853 14833 33891 14867
rect 33925 14833 33963 14867
rect 33997 14833 34035 14867
rect 34069 14833 34107 14867
rect 34141 14833 34179 14867
rect 34213 14833 34251 14867
rect 34285 14833 34323 14867
rect 34357 14833 34395 14867
rect 34429 14833 34467 14867
rect 34501 14833 34539 14867
rect 34573 14833 34611 14867
rect 34645 14833 34683 14867
rect 34717 14833 34755 14867
rect 34789 14833 34827 14867
rect 34861 14833 34899 14867
rect 34933 14833 34971 14867
rect 35005 14833 35043 14867
rect 35077 14833 35115 14867
rect 35149 14833 35187 14867
rect 35221 14833 35240 14867
rect -17320 14820 35240 14833
rect -17480 14797 -17420 14800
rect -17480 14763 -17467 14797
rect -17433 14763 -17420 14797
rect -17480 14725 -17420 14763
rect -17480 14691 -17467 14725
rect -17433 14691 -17420 14725
rect -17480 14653 -17420 14691
rect -17480 14619 -17467 14653
rect -17433 14619 -17420 14653
rect -17480 14581 -17420 14619
rect -17480 14547 -17467 14581
rect -17433 14547 -17420 14581
rect -17480 14509 -17420 14547
rect -17480 14475 -17467 14509
rect -17433 14475 -17420 14509
rect -17480 14437 -17420 14475
rect -17480 14403 -17467 14437
rect -17433 14403 -17420 14437
rect -17480 14365 -17420 14403
rect -17480 14331 -17467 14365
rect -17433 14331 -17420 14365
rect -17480 14293 -17420 14331
rect -17480 14259 -17467 14293
rect -17433 14259 -17420 14293
rect -17480 14221 -17420 14259
rect -17480 14187 -17467 14221
rect -17433 14187 -17420 14221
rect -17480 14149 -17420 14187
rect -17480 14115 -17467 14149
rect -17433 14115 -17420 14149
rect -17480 14077 -17420 14115
rect -17480 14043 -17467 14077
rect -17433 14043 -17420 14077
rect -17480 14005 -17420 14043
rect -17480 13971 -17467 14005
rect -17433 13971 -17420 14005
rect -17480 13933 -17420 13971
rect -17480 13920 -17467 13933
rect -17500 13899 -17467 13920
rect -17433 13920 -17420 13933
rect 35320 14797 35380 14800
rect 35320 14763 35333 14797
rect 35367 14763 35380 14797
rect 35320 14725 35380 14763
rect 35320 14691 35333 14725
rect 35367 14691 35380 14725
rect 35320 14653 35380 14691
rect 35320 14619 35333 14653
rect 35367 14619 35380 14653
rect 35320 14581 35380 14619
rect 35320 14547 35333 14581
rect 35367 14547 35380 14581
rect 35320 14509 35380 14547
rect 35320 14475 35333 14509
rect 35367 14475 35380 14509
rect 35320 14437 35380 14475
rect 35320 14403 35333 14437
rect 35367 14403 35380 14437
rect 35320 14365 35380 14403
rect 35320 14331 35333 14365
rect 35367 14331 35380 14365
rect 35320 14293 35380 14331
rect 35320 14259 35333 14293
rect 35367 14259 35380 14293
rect 35320 14221 35380 14259
rect 35320 14187 35333 14221
rect 35367 14187 35380 14221
rect 35320 14149 35380 14187
rect 35320 14115 35333 14149
rect 35367 14115 35380 14149
rect 35320 14077 35380 14115
rect 35320 14043 35333 14077
rect 35367 14043 35380 14077
rect 35320 14005 35380 14043
rect 35320 13971 35333 14005
rect 35367 13971 35380 14005
rect 35320 13933 35380 13971
rect 35320 13920 35333 13933
rect -17433 13899 35333 13920
rect 35367 13899 35380 13933
rect -17500 13861 35380 13899
rect -17500 13860 -17467 13861
rect -17480 13827 -17467 13860
rect -17433 13860 35333 13861
rect -17433 13827 -17420 13860
rect -17480 13789 -17420 13827
rect -17480 13755 -17467 13789
rect -17433 13755 -17420 13789
rect -17480 13717 -17420 13755
rect -17480 13683 -17467 13717
rect -17433 13683 -17420 13717
rect -17480 13645 -17420 13683
rect -17480 13611 -17467 13645
rect -17433 13611 -17420 13645
rect -17480 13573 -17420 13611
rect -17480 13539 -17467 13573
rect -17433 13539 -17420 13573
rect -17480 13501 -17420 13539
rect -17480 13467 -17467 13501
rect -17433 13467 -17420 13501
rect -17480 13429 -17420 13467
rect -17480 13395 -17467 13429
rect -17433 13395 -17420 13429
rect -17480 13357 -17420 13395
rect -17480 13323 -17467 13357
rect -17433 13323 -17420 13357
rect -17480 13285 -17420 13323
rect -17480 13251 -17467 13285
rect -17433 13251 -17420 13285
rect -17480 13213 -17420 13251
rect -17480 13179 -17467 13213
rect -17433 13179 -17420 13213
rect -17480 13141 -17420 13179
rect -17480 13107 -17467 13141
rect -17433 13107 -17420 13141
rect -17480 13069 -17420 13107
rect -17480 13035 -17467 13069
rect -17433 13035 -17420 13069
rect -17480 12997 -17420 13035
rect -17480 12963 -17467 12997
rect -17433 12963 -17420 12997
rect -17480 12925 -17420 12963
rect -17480 12891 -17467 12925
rect -17433 12891 -17420 12925
rect -17480 12853 -17420 12891
rect -17480 12819 -17467 12853
rect -17433 12819 -17420 12853
rect -17480 12781 -17420 12819
rect -17480 12747 -17467 12781
rect -17433 12747 -17420 12781
rect -17480 12709 -17420 12747
rect -17480 12675 -17467 12709
rect -17433 12675 -17420 12709
rect -17480 12637 -17420 12675
rect -17480 12603 -17467 12637
rect -17433 12603 -17420 12637
rect -17480 12565 -17420 12603
rect -17480 12531 -17467 12565
rect -17433 12531 -17420 12565
rect -17480 12493 -17420 12531
rect -17480 12459 -17467 12493
rect -17433 12459 -17420 12493
rect -17480 12421 -17420 12459
rect -17480 12387 -17467 12421
rect -17433 12387 -17420 12421
rect -17480 12349 -17420 12387
rect -17480 12315 -17467 12349
rect -17433 12315 -17420 12349
rect -17480 12277 -17420 12315
rect -17480 12243 -17467 12277
rect -17433 12243 -17420 12277
rect -17480 12205 -17420 12243
rect -17480 12171 -17467 12205
rect -17433 12171 -17420 12205
rect -17480 12133 -17420 12171
rect -17480 12100 -17467 12133
rect -17500 12099 -17467 12100
rect -17433 12100 -17420 12133
rect 35320 13827 35333 13860
rect 35367 13827 35380 13861
rect 35320 13789 35380 13827
rect 35320 13755 35333 13789
rect 35367 13755 35380 13789
rect 35320 13717 35380 13755
rect 35320 13683 35333 13717
rect 35367 13683 35380 13717
rect 35320 13645 35380 13683
rect 35320 13611 35333 13645
rect 35367 13611 35380 13645
rect 35320 13573 35380 13611
rect 35320 13539 35333 13573
rect 35367 13539 35380 13573
rect 35320 13501 35380 13539
rect 35320 13467 35333 13501
rect 35367 13467 35380 13501
rect 35320 13429 35380 13467
rect 35320 13395 35333 13429
rect 35367 13395 35380 13429
rect 35320 13357 35380 13395
rect 35320 13323 35333 13357
rect 35367 13323 35380 13357
rect 35320 13285 35380 13323
rect 35320 13251 35333 13285
rect 35367 13251 35380 13285
rect 35320 13213 35380 13251
rect 35320 13179 35333 13213
rect 35367 13179 35380 13213
rect 35320 13141 35380 13179
rect 35320 13107 35333 13141
rect 35367 13107 35380 13141
rect 35320 13069 35380 13107
rect 35320 13035 35333 13069
rect 35367 13035 35380 13069
rect 35320 12997 35380 13035
rect 35320 12963 35333 12997
rect 35367 12963 35380 12997
rect 35320 12925 35380 12963
rect 35320 12891 35333 12925
rect 35367 12891 35380 12925
rect 35320 12853 35380 12891
rect 35320 12819 35333 12853
rect 35367 12819 35380 12853
rect 35320 12781 35380 12819
rect 35320 12747 35333 12781
rect 35367 12747 35380 12781
rect 35320 12709 35380 12747
rect 35320 12675 35333 12709
rect 35367 12675 35380 12709
rect 35320 12637 35380 12675
rect 35320 12603 35333 12637
rect 35367 12603 35380 12637
rect 35320 12565 35380 12603
rect 35320 12531 35333 12565
rect 35367 12531 35380 12565
rect 35320 12493 35380 12531
rect 35320 12459 35333 12493
rect 35367 12459 35380 12493
rect 35320 12421 35380 12459
rect 35320 12387 35333 12421
rect 35367 12387 35380 12421
rect 35320 12349 35380 12387
rect 35320 12315 35333 12349
rect 35367 12315 35380 12349
rect 35320 12277 35380 12315
rect 35320 12243 35333 12277
rect 35367 12243 35380 12277
rect 35320 12205 35380 12243
rect 35320 12171 35333 12205
rect 35367 12171 35380 12205
rect 35320 12133 35380 12171
rect 35320 12100 35333 12133
rect -17433 12099 35333 12100
rect 35367 12100 35380 12133
rect 35367 12099 35400 12100
rect -17500 12061 35400 12099
rect -17500 12040 -17467 12061
rect -17480 12027 -17467 12040
rect -17433 12040 35333 12061
rect -17433 12027 -17420 12040
rect -17480 11989 -17420 12027
rect -17480 11955 -17467 11989
rect -17433 11955 -17420 11989
rect -17480 11917 -17420 11955
rect -17480 11883 -17467 11917
rect -17433 11883 -17420 11917
rect -17480 11845 -17420 11883
rect -17480 11811 -17467 11845
rect -17433 11811 -17420 11845
rect -17480 11773 -17420 11811
rect -17480 11739 -17467 11773
rect -17433 11739 -17420 11773
rect -17480 11701 -17420 11739
rect -17480 11667 -17467 11701
rect -17433 11667 -17420 11701
rect -17480 11629 -17420 11667
rect -17480 11595 -17467 11629
rect -17433 11595 -17420 11629
rect -17480 11557 -17420 11595
rect -17480 11523 -17467 11557
rect -17433 11523 -17420 11557
rect -17480 11485 -17420 11523
rect -17480 11451 -17467 11485
rect -17433 11451 -17420 11485
rect -17480 11413 -17420 11451
rect -17480 11379 -17467 11413
rect -17433 11379 -17420 11413
rect -17480 11341 -17420 11379
rect -17480 11307 -17467 11341
rect -17433 11307 -17420 11341
rect -17480 11269 -17420 11307
rect -17480 11235 -17467 11269
rect -17433 11235 -17420 11269
rect -17480 11197 -17420 11235
rect -17480 11163 -17467 11197
rect -17433 11163 -17420 11197
rect -17480 11125 -17420 11163
rect -17480 11091 -17467 11125
rect -17433 11091 -17420 11125
rect -17480 11053 -17420 11091
rect -17480 11019 -17467 11053
rect -17433 11019 -17420 11053
rect -17480 10981 -17420 11019
rect -17480 10947 -17467 10981
rect -17433 10947 -17420 10981
rect -17480 10909 -17420 10947
rect -17480 10875 -17467 10909
rect -17433 10875 -17420 10909
rect -17480 10837 -17420 10875
rect -17480 10803 -17467 10837
rect -17433 10803 -17420 10837
rect -17480 10765 -17420 10803
rect -17480 10731 -17467 10765
rect -17433 10731 -17420 10765
rect -17480 10693 -17420 10731
rect -17480 10659 -17467 10693
rect -17433 10659 -17420 10693
rect -17480 10621 -17420 10659
rect -17480 10587 -17467 10621
rect -17433 10587 -17420 10621
rect -17480 10549 -17420 10587
rect -17480 10515 -17467 10549
rect -17433 10515 -17420 10549
rect -17480 10477 -17420 10515
rect -17480 10443 -17467 10477
rect -17433 10443 -17420 10477
rect -17480 10420 -17420 10443
rect 35320 12027 35333 12040
rect 35367 12040 35400 12061
rect 35367 12027 35380 12040
rect 35320 11989 35380 12027
rect 35320 11955 35333 11989
rect 35367 11955 35380 11989
rect 35320 11917 35380 11955
rect 35320 11883 35333 11917
rect 35367 11883 35380 11917
rect 35320 11845 35380 11883
rect 35320 11811 35333 11845
rect 35367 11811 35380 11845
rect 35320 11773 35380 11811
rect 35320 11739 35333 11773
rect 35367 11739 35380 11773
rect 35320 11701 35380 11739
rect 35320 11667 35333 11701
rect 35367 11667 35380 11701
rect 35320 11629 35380 11667
rect 35320 11595 35333 11629
rect 35367 11595 35380 11629
rect 35320 11557 35380 11595
rect 35320 11523 35333 11557
rect 35367 11523 35380 11557
rect 35320 11485 35380 11523
rect 35320 11451 35333 11485
rect 35367 11451 35380 11485
rect 35320 11413 35380 11451
rect 35320 11379 35333 11413
rect 35367 11379 35380 11413
rect 35320 11341 35380 11379
rect 35320 11307 35333 11341
rect 35367 11307 35380 11341
rect 35320 11269 35380 11307
rect 35320 11235 35333 11269
rect 35367 11235 35380 11269
rect 35320 11197 35380 11235
rect 35320 11163 35333 11197
rect 35367 11163 35380 11197
rect 35320 11125 35380 11163
rect 35320 11091 35333 11125
rect 35367 11091 35380 11125
rect 35320 11053 35380 11091
rect 35320 11019 35333 11053
rect 35367 11019 35380 11053
rect 35320 10981 35380 11019
rect 35320 10947 35333 10981
rect 35367 10947 35380 10981
rect 35320 10909 35380 10947
rect 35320 10875 35333 10909
rect 35367 10875 35380 10909
rect 35320 10837 35380 10875
rect 35320 10803 35333 10837
rect 35367 10803 35380 10837
rect 35320 10765 35380 10803
rect 35320 10731 35333 10765
rect 35367 10731 35380 10765
rect 35320 10693 35380 10731
rect 35320 10659 35333 10693
rect 35367 10659 35380 10693
rect 35320 10621 35380 10659
rect 35320 10587 35333 10621
rect 35367 10587 35380 10621
rect 35320 10549 35380 10587
rect 35320 10515 35333 10549
rect 35367 10515 35380 10549
rect 35320 10477 35380 10515
rect 35320 10443 35333 10477
rect 35367 10443 35380 10477
rect 35320 10420 35380 10443
rect -17500 10405 35400 10420
rect -17500 10371 -17467 10405
rect -17433 10371 35333 10405
rect 35367 10371 35400 10405
rect -17500 10360 35400 10371
rect -17480 10333 -17420 10360
rect -17480 10299 -17467 10333
rect -17433 10299 -17420 10333
rect -17480 10261 -17420 10299
rect -17480 10227 -17467 10261
rect -17433 10227 -17420 10261
rect -17480 10189 -17420 10227
rect -17480 10155 -17467 10189
rect -17433 10155 -17420 10189
rect -17480 10117 -17420 10155
rect -17480 10083 -17467 10117
rect -17433 10083 -17420 10117
rect -17480 10045 -17420 10083
rect -17480 10011 -17467 10045
rect -17433 10011 -17420 10045
rect -17480 9973 -17420 10011
rect -17480 9939 -17467 9973
rect -17433 9939 -17420 9973
rect -17480 9901 -17420 9939
rect -17480 9867 -17467 9901
rect -17433 9867 -17420 9901
rect -17480 9829 -17420 9867
rect -17480 9795 -17467 9829
rect -17433 9795 -17420 9829
rect -17480 9757 -17420 9795
rect -17480 9723 -17467 9757
rect -17433 9723 -17420 9757
rect -17480 9685 -17420 9723
rect -17480 9651 -17467 9685
rect -17433 9651 -17420 9685
rect -17480 9613 -17420 9651
rect -17480 9579 -17467 9613
rect -17433 9579 -17420 9613
rect -17480 9541 -17420 9579
rect -17480 9507 -17467 9541
rect -17433 9507 -17420 9541
rect -17480 9469 -17420 9507
rect -17480 9435 -17467 9469
rect -17433 9435 -17420 9469
rect -17480 9397 -17420 9435
rect -17480 9363 -17467 9397
rect -17433 9363 -17420 9397
rect -17480 9325 -17420 9363
rect -17480 9291 -17467 9325
rect -17433 9291 -17420 9325
rect -17480 9253 -17420 9291
rect -17480 9219 -17467 9253
rect -17433 9219 -17420 9253
rect -17480 9181 -17420 9219
rect -17480 9147 -17467 9181
rect -17433 9147 -17420 9181
rect -17480 9109 -17420 9147
rect -17480 9075 -17467 9109
rect -17433 9075 -17420 9109
rect -17480 9037 -17420 9075
rect -17480 9003 -17467 9037
rect -17433 9003 -17420 9037
rect -17480 8965 -17420 9003
rect -17480 8931 -17467 8965
rect -17433 8931 -17420 8965
rect -17480 8893 -17420 8931
rect -17480 8859 -17467 8893
rect -17433 8859 -17420 8893
rect -17480 8821 -17420 8859
rect -17480 8787 -17467 8821
rect -17433 8787 -17420 8821
rect -17480 8749 -17420 8787
rect -17480 8715 -17467 8749
rect -17433 8715 -17420 8749
rect -17480 8677 -17420 8715
rect -17480 8643 -17467 8677
rect -17433 8643 -17420 8677
rect -17480 8605 -17420 8643
rect -17480 8600 -17467 8605
rect -17500 8571 -17467 8600
rect -17433 8600 -17420 8605
rect 35320 10333 35380 10360
rect 35320 10299 35333 10333
rect 35367 10299 35380 10333
rect 35320 10261 35380 10299
rect 35320 10227 35333 10261
rect 35367 10227 35380 10261
rect 35320 10189 35380 10227
rect 35320 10155 35333 10189
rect 35367 10155 35380 10189
rect 35320 10117 35380 10155
rect 35320 10083 35333 10117
rect 35367 10083 35380 10117
rect 35320 10045 35380 10083
rect 35320 10011 35333 10045
rect 35367 10011 35380 10045
rect 35320 9973 35380 10011
rect 35320 9939 35333 9973
rect 35367 9939 35380 9973
rect 35320 9901 35380 9939
rect 35320 9867 35333 9901
rect 35367 9867 35380 9901
rect 35320 9829 35380 9867
rect 35320 9795 35333 9829
rect 35367 9795 35380 9829
rect 35320 9757 35380 9795
rect 35320 9723 35333 9757
rect 35367 9723 35380 9757
rect 35320 9685 35380 9723
rect 35320 9651 35333 9685
rect 35367 9651 35380 9685
rect 35320 9613 35380 9651
rect 35320 9579 35333 9613
rect 35367 9579 35380 9613
rect 35320 9541 35380 9579
rect 35320 9507 35333 9541
rect 35367 9507 35380 9541
rect 35320 9469 35380 9507
rect 35320 9435 35333 9469
rect 35367 9435 35380 9469
rect 35320 9397 35380 9435
rect 35320 9363 35333 9397
rect 35367 9363 35380 9397
rect 35320 9325 35380 9363
rect 35320 9291 35333 9325
rect 35367 9291 35380 9325
rect 35320 9253 35380 9291
rect 35320 9219 35333 9253
rect 35367 9219 35380 9253
rect 35320 9181 35380 9219
rect 35320 9147 35333 9181
rect 35367 9147 35380 9181
rect 35320 9109 35380 9147
rect 35320 9075 35333 9109
rect 35367 9075 35380 9109
rect 35320 9037 35380 9075
rect 35320 9003 35333 9037
rect 35367 9003 35380 9037
rect 35320 8965 35380 9003
rect 35320 8931 35333 8965
rect 35367 8931 35380 8965
rect 35320 8893 35380 8931
rect 35320 8859 35333 8893
rect 35367 8859 35380 8893
rect 35320 8821 35380 8859
rect 35320 8787 35333 8821
rect 35367 8787 35380 8821
rect 35320 8749 35380 8787
rect 35320 8715 35333 8749
rect 35367 8715 35380 8749
rect 35320 8677 35380 8715
rect 35320 8643 35333 8677
rect 35367 8643 35380 8677
rect 35320 8605 35380 8643
rect 35320 8600 35333 8605
rect -17433 8571 35333 8600
rect 35367 8600 35380 8605
rect 35367 8571 35400 8600
rect -17500 8540 35400 8571
rect -17480 8533 -17420 8540
rect -17480 8499 -17467 8533
rect -17433 8499 -17420 8533
rect -17480 8461 -17420 8499
rect -17480 8427 -17467 8461
rect -17433 8427 -17420 8461
rect -17480 8389 -17420 8427
rect -17480 8355 -17467 8389
rect -17433 8355 -17420 8389
rect -17480 8317 -17420 8355
rect -17480 8283 -17467 8317
rect -17433 8283 -17420 8317
rect -17480 8245 -17420 8283
rect -17480 8211 -17467 8245
rect -17433 8211 -17420 8245
rect -17480 8173 -17420 8211
rect -17480 8139 -17467 8173
rect -17433 8139 -17420 8173
rect -17480 8101 -17420 8139
rect -17480 8067 -17467 8101
rect -17433 8067 -17420 8101
rect -17480 8029 -17420 8067
rect -17480 7995 -17467 8029
rect -17433 7995 -17420 8029
rect -17480 7957 -17420 7995
rect -17480 7923 -17467 7957
rect -17433 7923 -17420 7957
rect -17480 7885 -17420 7923
rect -17480 7851 -17467 7885
rect -17433 7851 -17420 7885
rect -17480 7813 -17420 7851
rect -17480 7779 -17467 7813
rect -17433 7779 -17420 7813
rect -17480 7741 -17420 7779
rect -17480 7707 -17467 7741
rect -17433 7707 -17420 7741
rect -17480 7669 -17420 7707
rect -17480 7635 -17467 7669
rect -17433 7635 -17420 7669
rect -17480 7597 -17420 7635
rect -17480 7563 -17467 7597
rect -17433 7563 -17420 7597
rect -17480 7525 -17420 7563
rect -17480 7491 -17467 7525
rect -17433 7491 -17420 7525
rect -17480 7453 -17420 7491
rect -17480 7419 -17467 7453
rect -17433 7419 -17420 7453
rect -17480 7381 -17420 7419
rect -17480 7347 -17467 7381
rect -17433 7347 -17420 7381
rect -17480 7309 -17420 7347
rect -17480 7275 -17467 7309
rect -17433 7275 -17420 7309
rect -17480 7237 -17420 7275
rect -17480 7203 -17467 7237
rect -17433 7203 -17420 7237
rect -17480 7165 -17420 7203
rect -17480 7131 -17467 7165
rect -17433 7131 -17420 7165
rect -17480 7093 -17420 7131
rect -17480 7059 -17467 7093
rect -17433 7059 -17420 7093
rect -17480 7021 -17420 7059
rect -17480 6987 -17467 7021
rect -17433 6987 -17420 7021
rect -17480 6949 -17420 6987
rect -17480 6915 -17467 6949
rect -17433 6915 -17420 6949
rect -17480 6877 -17420 6915
rect -17480 6843 -17467 6877
rect -17433 6843 -17420 6877
rect -17480 6805 -17420 6843
rect -17480 6771 -17467 6805
rect -17433 6771 -17420 6805
rect -17480 6733 -17420 6771
rect -17480 6699 -17467 6733
rect -17433 6699 -17420 6733
rect -17480 6661 -17420 6699
rect -17480 6627 -17467 6661
rect -17433 6627 -17420 6661
rect -17480 6589 -17420 6627
rect -17480 6555 -17467 6589
rect -17433 6555 -17420 6589
rect -17480 6520 -17420 6555
rect 35320 8533 35380 8540
rect 35320 8499 35333 8533
rect 35367 8499 35380 8533
rect 35320 8461 35380 8499
rect 35320 8427 35333 8461
rect 35367 8427 35380 8461
rect 35320 8389 35380 8427
rect 35320 8355 35333 8389
rect 35367 8355 35380 8389
rect 35320 8317 35380 8355
rect 35320 8283 35333 8317
rect 35367 8283 35380 8317
rect 35320 8245 35380 8283
rect 35320 8211 35333 8245
rect 35367 8211 35380 8245
rect 35320 8173 35380 8211
rect 35320 8139 35333 8173
rect 35367 8139 35380 8173
rect 35320 8101 35380 8139
rect 35320 8067 35333 8101
rect 35367 8067 35380 8101
rect 35320 8029 35380 8067
rect 35320 7995 35333 8029
rect 35367 7995 35380 8029
rect 35320 7957 35380 7995
rect 35320 7923 35333 7957
rect 35367 7923 35380 7957
rect 35320 7885 35380 7923
rect 35320 7851 35333 7885
rect 35367 7851 35380 7885
rect 35320 7813 35380 7851
rect 35320 7779 35333 7813
rect 35367 7779 35380 7813
rect 35320 7741 35380 7779
rect 35320 7707 35333 7741
rect 35367 7707 35380 7741
rect 35320 7669 35380 7707
rect 35320 7635 35333 7669
rect 35367 7635 35380 7669
rect 35320 7597 35380 7635
rect 35320 7563 35333 7597
rect 35367 7563 35380 7597
rect 35320 7525 35380 7563
rect 35320 7491 35333 7525
rect 35367 7491 35380 7525
rect 35320 7453 35380 7491
rect 35320 7419 35333 7453
rect 35367 7419 35380 7453
rect 35320 7381 35380 7419
rect 35320 7347 35333 7381
rect 35367 7347 35380 7381
rect 35320 7309 35380 7347
rect 35320 7275 35333 7309
rect 35367 7275 35380 7309
rect 35320 7237 35380 7275
rect 35320 7203 35333 7237
rect 35367 7203 35380 7237
rect 35320 7165 35380 7203
rect 35320 7131 35333 7165
rect 35367 7131 35380 7165
rect 35320 7093 35380 7131
rect 35320 7059 35333 7093
rect 35367 7059 35380 7093
rect 35320 7021 35380 7059
rect 35320 6987 35333 7021
rect 35367 6987 35380 7021
rect 35320 6949 35380 6987
rect 35320 6915 35333 6949
rect 35367 6915 35380 6949
rect 35320 6877 35380 6915
rect 35320 6843 35333 6877
rect 35367 6843 35380 6877
rect 35320 6805 35380 6843
rect 35320 6771 35333 6805
rect 35367 6771 35380 6805
rect 35320 6733 35380 6771
rect 35320 6699 35333 6733
rect 35367 6699 35380 6733
rect 35320 6661 35380 6699
rect 35320 6627 35333 6661
rect 35367 6627 35380 6661
rect 35320 6589 35380 6627
rect 35320 6555 35333 6589
rect 35367 6555 35380 6589
rect 35320 6520 35380 6555
rect -17500 6517 200 6520
rect -17500 6483 -17467 6517
rect -17433 6483 200 6517
rect -17500 6460 200 6483
rect 17700 6517 35400 6520
rect 17700 6483 35333 6517
rect 35367 6483 35400 6517
rect 17700 6460 35400 6483
rect -17480 6445 -17420 6460
rect -17480 6411 -17467 6445
rect -17433 6411 -17420 6445
rect -17480 6373 -17420 6411
rect -17480 6339 -17467 6373
rect -17433 6339 -17420 6373
rect -17480 6301 -17420 6339
rect -17480 6267 -17467 6301
rect -17433 6267 -17420 6301
rect -17480 6229 -17420 6267
rect -17480 6195 -17467 6229
rect -17433 6195 -17420 6229
rect -17480 6157 -17420 6195
rect -17480 6123 -17467 6157
rect -17433 6123 -17420 6157
rect -17480 6085 -17420 6123
rect -17480 6051 -17467 6085
rect -17433 6051 -17420 6085
rect -17480 6013 -17420 6051
rect -17480 5979 -17467 6013
rect -17433 5979 -17420 6013
rect -17480 5941 -17420 5979
rect -17480 5907 -17467 5941
rect -17433 5907 -17420 5941
rect -17480 5869 -17420 5907
rect -17480 5835 -17467 5869
rect -17433 5835 -17420 5869
rect -17480 5797 -17420 5835
rect -17480 5763 -17467 5797
rect -17433 5763 -17420 5797
rect -17480 5725 -17420 5763
rect -17480 5691 -17467 5725
rect -17433 5691 -17420 5725
rect -17480 5653 -17420 5691
rect -17480 5619 -17467 5653
rect -17433 5619 -17420 5653
rect -17480 5581 -17420 5619
rect -17480 5547 -17467 5581
rect -17433 5547 -17420 5581
rect -17480 5509 -17420 5547
rect -17480 5475 -17467 5509
rect -17433 5475 -17420 5509
rect -17480 5437 -17420 5475
rect -17480 5403 -17467 5437
rect -17433 5403 -17420 5437
rect -17480 5365 -17420 5403
rect -17480 5331 -17467 5365
rect -17433 5331 -17420 5365
rect -17480 5293 -17420 5331
rect -17480 5259 -17467 5293
rect -17433 5259 -17420 5293
rect -17480 5221 -17420 5259
rect -17480 5187 -17467 5221
rect -17433 5187 -17420 5221
rect -17480 5149 -17420 5187
rect -17480 5115 -17467 5149
rect -17433 5115 -17420 5149
rect -17480 5077 -17420 5115
rect -17480 5043 -17467 5077
rect -17433 5043 -17420 5077
rect -17480 5005 -17420 5043
rect -17480 4971 -17467 5005
rect -17433 4971 -17420 5005
rect -17480 4933 -17420 4971
rect -17480 4899 -17467 4933
rect -17433 4899 -17420 4933
rect -17480 4861 -17420 4899
rect -17480 4827 -17467 4861
rect -17433 4827 -17420 4861
rect -17480 4789 -17420 4827
rect -17480 4755 -17467 4789
rect -17433 4755 -17420 4789
rect -17480 4717 -17420 4755
rect -17480 4700 -17467 4717
rect -17500 4683 -17467 4700
rect -17433 4700 -17420 4717
rect 35320 6445 35380 6460
rect 35320 6411 35333 6445
rect 35367 6411 35380 6445
rect 35320 6373 35380 6411
rect 35320 6339 35333 6373
rect 35367 6339 35380 6373
rect 35320 6301 35380 6339
rect 35320 6267 35333 6301
rect 35367 6267 35380 6301
rect 35320 6229 35380 6267
rect 35320 6195 35333 6229
rect 35367 6195 35380 6229
rect 35320 6157 35380 6195
rect 35320 6123 35333 6157
rect 35367 6123 35380 6157
rect 35320 6085 35380 6123
rect 35320 6051 35333 6085
rect 35367 6051 35380 6085
rect 35320 6013 35380 6051
rect 35320 5979 35333 6013
rect 35367 5979 35380 6013
rect 35320 5941 35380 5979
rect 35320 5907 35333 5941
rect 35367 5907 35380 5941
rect 35320 5869 35380 5907
rect 35320 5835 35333 5869
rect 35367 5835 35380 5869
rect 35320 5797 35380 5835
rect 35320 5763 35333 5797
rect 35367 5763 35380 5797
rect 35320 5725 35380 5763
rect 35320 5691 35333 5725
rect 35367 5691 35380 5725
rect 35320 5653 35380 5691
rect 35320 5619 35333 5653
rect 35367 5619 35380 5653
rect 35320 5581 35380 5619
rect 35320 5547 35333 5581
rect 35367 5547 35380 5581
rect 35320 5509 35380 5547
rect 35320 5475 35333 5509
rect 35367 5475 35380 5509
rect 35320 5437 35380 5475
rect 35320 5403 35333 5437
rect 35367 5403 35380 5437
rect 35320 5365 35380 5403
rect 35320 5331 35333 5365
rect 35367 5331 35380 5365
rect 35320 5293 35380 5331
rect 35320 5259 35333 5293
rect 35367 5259 35380 5293
rect 35320 5221 35380 5259
rect 35320 5187 35333 5221
rect 35367 5187 35380 5221
rect 35320 5149 35380 5187
rect 35320 5115 35333 5149
rect 35367 5115 35380 5149
rect 35320 5077 35380 5115
rect 35320 5043 35333 5077
rect 35367 5043 35380 5077
rect 35320 5005 35380 5043
rect 35320 4971 35333 5005
rect 35367 4971 35380 5005
rect 35320 4933 35380 4971
rect 35320 4899 35333 4933
rect 35367 4899 35380 4933
rect 35320 4861 35380 4899
rect 35320 4827 35333 4861
rect 35367 4827 35380 4861
rect 35320 4789 35380 4827
rect 35320 4755 35333 4789
rect 35367 4755 35380 4789
rect 35320 4717 35380 4755
rect 35320 4700 35333 4717
rect -17433 4683 200 4700
rect -17500 4645 200 4683
rect -17500 4640 -17467 4645
rect -17480 4611 -17467 4640
rect -17433 4640 200 4645
rect 17700 4683 35333 4700
rect 35367 4700 35380 4717
rect 35367 4683 35400 4700
rect 17700 4645 35400 4683
rect 17700 4640 35333 4645
rect -17433 4611 -17420 4640
rect -17480 4573 -17420 4611
rect -17480 4539 -17467 4573
rect -17433 4539 -17420 4573
rect -17480 4501 -17420 4539
rect -17480 4467 -17467 4501
rect -17433 4467 -17420 4501
rect -17480 4429 -17420 4467
rect -17480 4395 -17467 4429
rect -17433 4395 -17420 4429
rect -17480 4357 -17420 4395
rect -17480 4323 -17467 4357
rect -17433 4323 -17420 4357
rect -17480 4285 -17420 4323
rect -17480 4251 -17467 4285
rect -17433 4251 -17420 4285
rect -17480 4213 -17420 4251
rect -17480 4179 -17467 4213
rect -17433 4179 -17420 4213
rect -17480 4141 -17420 4179
rect -17480 4107 -17467 4141
rect -17433 4107 -17420 4141
rect -17480 4069 -17420 4107
rect -17480 4035 -17467 4069
rect -17433 4035 -17420 4069
rect -17480 3997 -17420 4035
rect -17480 3963 -17467 3997
rect -17433 3963 -17420 3997
rect -17480 3925 -17420 3963
rect -17480 3891 -17467 3925
rect -17433 3891 -17420 3925
rect -17480 3853 -17420 3891
rect -17480 3819 -17467 3853
rect -17433 3819 -17420 3853
rect -17480 3781 -17420 3819
rect -17480 3747 -17467 3781
rect -17433 3747 -17420 3781
rect -17480 3709 -17420 3747
rect -17480 3675 -17467 3709
rect -17433 3675 -17420 3709
rect -17480 3637 -17420 3675
rect -17480 3603 -17467 3637
rect -17433 3603 -17420 3637
rect -17480 3565 -17420 3603
rect -17480 3531 -17467 3565
rect -17433 3531 -17420 3565
rect -17480 3493 -17420 3531
rect -17480 3459 -17467 3493
rect -17433 3459 -17420 3493
rect -17480 3421 -17420 3459
rect -17480 3387 -17467 3421
rect -17433 3387 -17420 3421
rect -17480 3349 -17420 3387
rect -17480 3315 -17467 3349
rect -17433 3315 -17420 3349
rect -17480 3277 -17420 3315
rect -17480 3243 -17467 3277
rect -17433 3243 -17420 3277
rect -17480 3205 -17420 3243
rect -17480 3171 -17467 3205
rect -17433 3171 -17420 3205
rect -17480 3133 -17420 3171
rect -17480 3099 -17467 3133
rect -17433 3099 -17420 3133
rect -17480 3061 -17420 3099
rect -17480 3027 -17467 3061
rect -17433 3027 -17420 3061
rect -17480 3020 -17420 3027
rect 35320 4611 35333 4640
rect 35367 4640 35400 4645
rect 35367 4611 35380 4640
rect 35320 4573 35380 4611
rect 35320 4539 35333 4573
rect 35367 4539 35380 4573
rect 35320 4501 35380 4539
rect 35320 4467 35333 4501
rect 35367 4467 35380 4501
rect 35320 4429 35380 4467
rect 35320 4395 35333 4429
rect 35367 4395 35380 4429
rect 35320 4357 35380 4395
rect 35320 4323 35333 4357
rect 35367 4323 35380 4357
rect 35320 4285 35380 4323
rect 35320 4251 35333 4285
rect 35367 4251 35380 4285
rect 35320 4213 35380 4251
rect 35320 4179 35333 4213
rect 35367 4179 35380 4213
rect 35320 4141 35380 4179
rect 35320 4107 35333 4141
rect 35367 4107 35380 4141
rect 35320 4069 35380 4107
rect 35320 4035 35333 4069
rect 35367 4035 35380 4069
rect 35320 3997 35380 4035
rect 35320 3963 35333 3997
rect 35367 3963 35380 3997
rect 35320 3925 35380 3963
rect 35320 3891 35333 3925
rect 35367 3891 35380 3925
rect 35320 3853 35380 3891
rect 35320 3819 35333 3853
rect 35367 3819 35380 3853
rect 35320 3781 35380 3819
rect 35320 3747 35333 3781
rect 35367 3747 35380 3781
rect 35320 3709 35380 3747
rect 35320 3675 35333 3709
rect 35367 3675 35380 3709
rect 35320 3637 35380 3675
rect 35320 3603 35333 3637
rect 35367 3603 35380 3637
rect 35320 3565 35380 3603
rect 35320 3531 35333 3565
rect 35367 3531 35380 3565
rect 35320 3493 35380 3531
rect 35320 3459 35333 3493
rect 35367 3459 35380 3493
rect 35320 3421 35380 3459
rect 35320 3387 35333 3421
rect 35367 3387 35380 3421
rect 35320 3349 35380 3387
rect 35320 3315 35333 3349
rect 35367 3315 35380 3349
rect 35320 3277 35380 3315
rect 35320 3243 35333 3277
rect 35367 3243 35380 3277
rect 35320 3205 35380 3243
rect 35320 3171 35333 3205
rect 35367 3171 35380 3205
rect 35320 3133 35380 3171
rect 35320 3099 35333 3133
rect 35367 3099 35380 3133
rect 35320 3061 35380 3099
rect 35320 3027 35333 3061
rect 35367 3027 35380 3061
rect 35320 3020 35380 3027
rect -17500 2989 200 3020
rect -17500 2960 -17467 2989
rect -17480 2955 -17467 2960
rect -17433 2960 200 2989
rect 17700 2989 35400 3020
rect 17700 2960 35333 2989
rect -17433 2955 -17420 2960
rect -17480 2917 -17420 2955
rect -17480 2883 -17467 2917
rect -17433 2883 -17420 2917
rect -17480 2845 -17420 2883
rect -17480 2811 -17467 2845
rect -17433 2811 -17420 2845
rect -17480 2773 -17420 2811
rect -17480 2739 -17467 2773
rect -17433 2739 -17420 2773
rect -17480 2701 -17420 2739
rect -17480 2667 -17467 2701
rect -17433 2667 -17420 2701
rect -17480 2629 -17420 2667
rect -17480 2595 -17467 2629
rect -17433 2595 -17420 2629
rect -17480 2557 -17420 2595
rect -17480 2523 -17467 2557
rect -17433 2523 -17420 2557
rect -17480 2485 -17420 2523
rect -17480 2451 -17467 2485
rect -17433 2451 -17420 2485
rect -17480 2413 -17420 2451
rect -17480 2379 -17467 2413
rect -17433 2379 -17420 2413
rect -17480 2341 -17420 2379
rect -17480 2307 -17467 2341
rect -17433 2307 -17420 2341
rect -17480 2269 -17420 2307
rect -17480 2235 -17467 2269
rect -17433 2235 -17420 2269
rect -17480 2197 -17420 2235
rect -17480 2163 -17467 2197
rect -17433 2163 -17420 2197
rect -17480 2125 -17420 2163
rect -17480 2091 -17467 2125
rect -17433 2091 -17420 2125
rect -17480 2053 -17420 2091
rect -17480 2019 -17467 2053
rect -17433 2019 -17420 2053
rect -17480 1981 -17420 2019
rect -17480 1947 -17467 1981
rect -17433 1947 -17420 1981
rect -17480 1909 -17420 1947
rect -17480 1875 -17467 1909
rect -17433 1875 -17420 1909
rect -17480 1837 -17420 1875
rect -17480 1803 -17467 1837
rect -17433 1803 -17420 1837
rect -17480 1765 -17420 1803
rect -17480 1731 -17467 1765
rect -17433 1731 -17420 1765
rect -17480 1693 -17420 1731
rect -17480 1659 -17467 1693
rect -17433 1659 -17420 1693
rect -17480 1621 -17420 1659
rect -17480 1587 -17467 1621
rect -17433 1587 -17420 1621
rect -17480 1549 -17420 1587
rect -17480 1515 -17467 1549
rect -17433 1515 -17420 1549
rect -17480 1477 -17420 1515
rect -17480 1443 -17467 1477
rect -17433 1443 -17420 1477
rect -17480 1405 -17420 1443
rect -17480 1371 -17467 1405
rect -17433 1371 -17420 1405
rect -17480 1333 -17420 1371
rect -17480 1299 -17467 1333
rect -17433 1299 -17420 1333
rect -17480 1261 -17420 1299
rect -17480 1227 -17467 1261
rect -17433 1227 -17420 1261
rect -17480 1200 -17420 1227
rect 35320 2955 35333 2960
rect 35367 2960 35400 2989
rect 35367 2955 35380 2960
rect 35320 2917 35380 2955
rect 35320 2883 35333 2917
rect 35367 2883 35380 2917
rect 35320 2845 35380 2883
rect 35320 2811 35333 2845
rect 35367 2811 35380 2845
rect 35320 2773 35380 2811
rect 35320 2739 35333 2773
rect 35367 2739 35380 2773
rect 35320 2701 35380 2739
rect 35320 2667 35333 2701
rect 35367 2667 35380 2701
rect 35320 2629 35380 2667
rect 35320 2595 35333 2629
rect 35367 2595 35380 2629
rect 35320 2557 35380 2595
rect 35320 2523 35333 2557
rect 35367 2523 35380 2557
rect 35320 2485 35380 2523
rect 35320 2451 35333 2485
rect 35367 2451 35380 2485
rect 35320 2413 35380 2451
rect 35320 2379 35333 2413
rect 35367 2379 35380 2413
rect 35320 2341 35380 2379
rect 35320 2307 35333 2341
rect 35367 2307 35380 2341
rect 35320 2269 35380 2307
rect 35320 2235 35333 2269
rect 35367 2235 35380 2269
rect 35320 2197 35380 2235
rect 35320 2163 35333 2197
rect 35367 2163 35380 2197
rect 35320 2125 35380 2163
rect 35320 2091 35333 2125
rect 35367 2091 35380 2125
rect 35320 2053 35380 2091
rect 35320 2019 35333 2053
rect 35367 2019 35380 2053
rect 35320 1981 35380 2019
rect 35320 1947 35333 1981
rect 35367 1947 35380 1981
rect 35320 1909 35380 1947
rect 35320 1875 35333 1909
rect 35367 1875 35380 1909
rect 35320 1837 35380 1875
rect 35320 1803 35333 1837
rect 35367 1803 35380 1837
rect 35320 1765 35380 1803
rect 35320 1731 35333 1765
rect 35367 1731 35380 1765
rect 35320 1693 35380 1731
rect 35320 1659 35333 1693
rect 35367 1659 35380 1693
rect 35320 1621 35380 1659
rect 35320 1587 35333 1621
rect 35367 1587 35380 1621
rect 35320 1549 35380 1587
rect 35320 1515 35333 1549
rect 35367 1515 35380 1549
rect 35320 1477 35380 1515
rect 35320 1443 35333 1477
rect 35367 1443 35380 1477
rect 35320 1405 35380 1443
rect 35320 1371 35333 1405
rect 35367 1371 35380 1405
rect 35320 1333 35380 1371
rect 35320 1299 35333 1333
rect 35367 1299 35380 1333
rect 35320 1261 35380 1299
rect 35320 1227 35333 1261
rect 35367 1227 35380 1261
rect 35320 1200 35380 1227
rect -17500 1189 200 1200
rect -17500 1155 -17467 1189
rect -17433 1155 200 1189
rect -17500 1140 200 1155
rect 17700 1189 35400 1200
rect 17700 1155 35333 1189
rect 35367 1155 35400 1189
rect 17700 1140 35400 1155
rect -17480 1117 -17420 1140
rect -17480 1083 -17467 1117
rect -17433 1083 -17420 1117
rect -17480 1045 -17420 1083
rect -17480 1011 -17467 1045
rect -17433 1011 -17420 1045
rect -17480 973 -17420 1011
rect -17480 939 -17467 973
rect -17433 939 -17420 973
rect -17480 901 -17420 939
rect -17480 867 -17467 901
rect -17433 867 -17420 901
rect -17480 829 -17420 867
rect -17480 795 -17467 829
rect -17433 795 -17420 829
rect -17480 757 -17420 795
rect -17480 723 -17467 757
rect -17433 723 -17420 757
rect -17480 685 -17420 723
rect -17480 651 -17467 685
rect -17433 651 -17420 685
rect -17480 613 -17420 651
rect -17480 579 -17467 613
rect -17433 579 -17420 613
rect -17480 541 -17420 579
rect -17480 507 -17467 541
rect -17433 507 -17420 541
rect -17480 469 -17420 507
rect -17480 435 -17467 469
rect -17433 435 -17420 469
rect -17480 397 -17420 435
rect -17480 363 -17467 397
rect -17433 363 -17420 397
rect -17480 325 -17420 363
rect -17480 291 -17467 325
rect -17433 291 -17420 325
rect -17480 253 -17420 291
rect -17480 219 -17467 253
rect -17433 219 -17420 253
rect -17480 181 -17420 219
rect -17480 147 -17467 181
rect -17433 147 -17420 181
rect -17480 109 -17420 147
rect -17480 75 -17467 109
rect -17433 75 -17420 109
rect -17480 37 -17420 75
rect -17480 3 -17467 37
rect -17433 3 -17420 37
rect -17480 -35 -17420 3
rect -17480 -69 -17467 -35
rect -17433 -69 -17420 -35
rect -17480 -107 -17420 -69
rect -17480 -141 -17467 -107
rect -17433 -141 -17420 -107
rect -17480 -179 -17420 -141
rect -17480 -213 -17467 -179
rect -17433 -213 -17420 -179
rect -17480 -251 -17420 -213
rect -17480 -285 -17467 -251
rect -17433 -285 -17420 -251
rect -17480 -323 -17420 -285
rect -17480 -357 -17467 -323
rect -17433 -357 -17420 -323
rect -17480 -395 -17420 -357
rect -17480 -429 -17467 -395
rect -17433 -429 -17420 -395
rect -17480 -467 -17420 -429
rect -17480 -501 -17467 -467
rect -17433 -501 -17420 -467
rect -17480 -539 -17420 -501
rect -17480 -573 -17467 -539
rect -17433 -573 -17420 -539
rect -17480 -611 -17420 -573
rect -17480 -645 -17467 -611
rect -17433 -645 -17420 -611
rect -17480 -683 -17420 -645
rect -17480 -717 -17467 -683
rect -17433 -717 -17420 -683
rect -17480 -755 -17420 -717
rect -17480 -789 -17467 -755
rect -17433 -789 -17420 -755
rect -17480 -827 -17420 -789
rect -17480 -861 -17467 -827
rect -17433 -861 -17420 -827
rect -17480 -880 -17420 -861
rect 35320 1117 35380 1140
rect 35320 1083 35333 1117
rect 35367 1083 35380 1117
rect 35320 1045 35380 1083
rect 35320 1011 35333 1045
rect 35367 1011 35380 1045
rect 35320 973 35380 1011
rect 35320 939 35333 973
rect 35367 939 35380 973
rect 35320 901 35380 939
rect 35320 867 35333 901
rect 35367 867 35380 901
rect 35320 829 35380 867
rect 35320 795 35333 829
rect 35367 795 35380 829
rect 35320 757 35380 795
rect 35320 723 35333 757
rect 35367 723 35380 757
rect 35320 685 35380 723
rect 35320 651 35333 685
rect 35367 651 35380 685
rect 35320 613 35380 651
rect 35320 579 35333 613
rect 35367 579 35380 613
rect 35320 541 35380 579
rect 35320 507 35333 541
rect 35367 507 35380 541
rect 35320 469 35380 507
rect 35320 435 35333 469
rect 35367 435 35380 469
rect 35320 397 35380 435
rect 35320 363 35333 397
rect 35367 363 35380 397
rect 35320 325 35380 363
rect 35320 291 35333 325
rect 35367 291 35380 325
rect 35320 253 35380 291
rect 35320 219 35333 253
rect 35367 219 35380 253
rect 35320 181 35380 219
rect 35320 147 35333 181
rect 35367 147 35380 181
rect 35320 109 35380 147
rect 35320 75 35333 109
rect 35367 75 35380 109
rect 35320 37 35380 75
rect 35320 3 35333 37
rect 35367 3 35380 37
rect 35320 -35 35380 3
rect 35320 -69 35333 -35
rect 35367 -69 35380 -35
rect 35320 -107 35380 -69
rect 35320 -141 35333 -107
rect 35367 -141 35380 -107
rect 35320 -179 35380 -141
rect 35320 -213 35333 -179
rect 35367 -213 35380 -179
rect 35320 -251 35380 -213
rect 35320 -285 35333 -251
rect 35367 -285 35380 -251
rect 35320 -323 35380 -285
rect 35320 -357 35333 -323
rect 35367 -357 35380 -323
rect 35320 -395 35380 -357
rect 35320 -429 35333 -395
rect 35367 -429 35380 -395
rect 35320 -467 35380 -429
rect 35320 -501 35333 -467
rect 35367 -501 35380 -467
rect 35320 -539 35380 -501
rect 35320 -573 35333 -539
rect 35367 -573 35380 -539
rect 35320 -611 35380 -573
rect 35320 -645 35333 -611
rect 35367 -645 35380 -611
rect 35320 -683 35380 -645
rect 35320 -717 35333 -683
rect 35367 -717 35380 -683
rect 35320 -755 35380 -717
rect 35320 -789 35333 -755
rect 35367 -789 35380 -755
rect 35320 -827 35380 -789
rect 35320 -861 35333 -827
rect 35367 -861 35380 -827
rect 35320 -880 35380 -861
rect -17500 -899 35400 -880
rect -17500 -933 -17467 -899
rect -17433 -933 35333 -899
rect 35367 -933 35400 -899
rect -17500 -940 35400 -933
rect -17480 -971 -17420 -940
rect -17480 -1005 -17467 -971
rect -17433 -1005 -17420 -971
rect -17480 -1043 -17420 -1005
rect -17480 -1077 -17467 -1043
rect -17433 -1077 -17420 -1043
rect -17480 -1115 -17420 -1077
rect -17480 -1149 -17467 -1115
rect -17433 -1149 -17420 -1115
rect -17480 -1187 -17420 -1149
rect -17480 -1221 -17467 -1187
rect -17433 -1221 -17420 -1187
rect -17480 -1259 -17420 -1221
rect -17480 -1293 -17467 -1259
rect -17433 -1293 -17420 -1259
rect -17480 -1331 -17420 -1293
rect -17480 -1365 -17467 -1331
rect -17433 -1365 -17420 -1331
rect -17480 -1403 -17420 -1365
rect -17480 -1437 -17467 -1403
rect -17433 -1437 -17420 -1403
rect -17480 -1475 -17420 -1437
rect -17480 -1509 -17467 -1475
rect -17433 -1509 -17420 -1475
rect -17480 -1547 -17420 -1509
rect -17480 -1581 -17467 -1547
rect -17433 -1581 -17420 -1547
rect -17480 -1619 -17420 -1581
rect -17480 -1653 -17467 -1619
rect -17433 -1653 -17420 -1619
rect -17480 -1691 -17420 -1653
rect -17480 -1725 -17467 -1691
rect -17433 -1725 -17420 -1691
rect -17480 -1763 -17420 -1725
rect -17480 -1797 -17467 -1763
rect -17433 -1797 -17420 -1763
rect -17480 -1835 -17420 -1797
rect -17480 -1869 -17467 -1835
rect -17433 -1869 -17420 -1835
rect -17480 -1907 -17420 -1869
rect -17480 -1941 -17467 -1907
rect -17433 -1941 -17420 -1907
rect -17480 -1979 -17420 -1941
rect -17480 -2013 -17467 -1979
rect -17433 -2013 -17420 -1979
rect -17480 -2051 -17420 -2013
rect -17480 -2085 -17467 -2051
rect -17433 -2085 -17420 -2051
rect -17480 -2123 -17420 -2085
rect -17480 -2157 -17467 -2123
rect -17433 -2157 -17420 -2123
rect -17480 -2195 -17420 -2157
rect -17480 -2229 -17467 -2195
rect -17433 -2229 -17420 -2195
rect -17480 -2267 -17420 -2229
rect -17480 -2301 -17467 -2267
rect -17433 -2301 -17420 -2267
rect -17480 -2339 -17420 -2301
rect -17480 -2373 -17467 -2339
rect -17433 -2373 -17420 -2339
rect -17480 -2411 -17420 -2373
rect -17480 -2445 -17467 -2411
rect -17433 -2445 -17420 -2411
rect -17480 -2483 -17420 -2445
rect -17480 -2517 -17467 -2483
rect -17433 -2517 -17420 -2483
rect -17480 -2555 -17420 -2517
rect -17480 -2589 -17467 -2555
rect -17433 -2589 -17420 -2555
rect -17480 -2627 -17420 -2589
rect -17480 -2661 -17467 -2627
rect -17433 -2661 -17420 -2627
rect -17480 -2699 -17420 -2661
rect -17480 -2700 -17467 -2699
rect -17500 -2733 -17467 -2700
rect -17433 -2700 -17420 -2699
rect 35320 -971 35380 -940
rect 35320 -1005 35333 -971
rect 35367 -1005 35380 -971
rect 35320 -1043 35380 -1005
rect 35320 -1077 35333 -1043
rect 35367 -1077 35380 -1043
rect 35320 -1115 35380 -1077
rect 35320 -1149 35333 -1115
rect 35367 -1149 35380 -1115
rect 35320 -1187 35380 -1149
rect 35320 -1221 35333 -1187
rect 35367 -1221 35380 -1187
rect 35320 -1259 35380 -1221
rect 35320 -1293 35333 -1259
rect 35367 -1293 35380 -1259
rect 35320 -1331 35380 -1293
rect 35320 -1365 35333 -1331
rect 35367 -1365 35380 -1331
rect 35320 -1403 35380 -1365
rect 35320 -1437 35333 -1403
rect 35367 -1437 35380 -1403
rect 35320 -1475 35380 -1437
rect 35320 -1509 35333 -1475
rect 35367 -1509 35380 -1475
rect 35320 -1547 35380 -1509
rect 35320 -1581 35333 -1547
rect 35367 -1581 35380 -1547
rect 35320 -1619 35380 -1581
rect 35320 -1653 35333 -1619
rect 35367 -1653 35380 -1619
rect 35320 -1691 35380 -1653
rect 35320 -1725 35333 -1691
rect 35367 -1725 35380 -1691
rect 35320 -1763 35380 -1725
rect 35320 -1797 35333 -1763
rect 35367 -1797 35380 -1763
rect 35320 -1835 35380 -1797
rect 35320 -1869 35333 -1835
rect 35367 -1869 35380 -1835
rect 35320 -1907 35380 -1869
rect 35320 -1941 35333 -1907
rect 35367 -1941 35380 -1907
rect 35320 -1979 35380 -1941
rect 35320 -2013 35333 -1979
rect 35367 -2013 35380 -1979
rect 35320 -2051 35380 -2013
rect 35320 -2085 35333 -2051
rect 35367 -2085 35380 -2051
rect 35320 -2123 35380 -2085
rect 35320 -2157 35333 -2123
rect 35367 -2157 35380 -2123
rect 35320 -2195 35380 -2157
rect 35320 -2229 35333 -2195
rect 35367 -2229 35380 -2195
rect 35320 -2267 35380 -2229
rect 35320 -2301 35333 -2267
rect 35367 -2301 35380 -2267
rect 35320 -2339 35380 -2301
rect 35320 -2373 35333 -2339
rect 35367 -2373 35380 -2339
rect 35320 -2411 35380 -2373
rect 35320 -2445 35333 -2411
rect 35367 -2445 35380 -2411
rect 35320 -2483 35380 -2445
rect 35320 -2517 35333 -2483
rect 35367 -2517 35380 -2483
rect 35320 -2555 35380 -2517
rect 35320 -2589 35333 -2555
rect 35367 -2589 35380 -2555
rect 35320 -2627 35380 -2589
rect 35320 -2661 35333 -2627
rect 35367 -2661 35380 -2627
rect 35320 -2699 35380 -2661
rect 35320 -2700 35333 -2699
rect -17433 -2733 35333 -2700
rect 35367 -2700 35380 -2699
rect 35367 -2733 35400 -2700
rect -17500 -2760 35400 -2733
rect -17480 -2771 -17420 -2760
rect -17480 -2805 -17467 -2771
rect -17433 -2805 -17420 -2771
rect -17480 -2843 -17420 -2805
rect -17480 -2877 -17467 -2843
rect -17433 -2877 -17420 -2843
rect -17480 -2915 -17420 -2877
rect -17480 -2949 -17467 -2915
rect -17433 -2949 -17420 -2915
rect -17480 -2987 -17420 -2949
rect -17480 -3021 -17467 -2987
rect -17433 -3021 -17420 -2987
rect -17480 -3059 -17420 -3021
rect -17480 -3093 -17467 -3059
rect -17433 -3093 -17420 -3059
rect -17480 -3131 -17420 -3093
rect -17480 -3165 -17467 -3131
rect -17433 -3165 -17420 -3131
rect -17480 -3203 -17420 -3165
rect -17480 -3237 -17467 -3203
rect -17433 -3237 -17420 -3203
rect -17480 -3275 -17420 -3237
rect -17480 -3309 -17467 -3275
rect -17433 -3309 -17420 -3275
rect -17480 -3347 -17420 -3309
rect -17480 -3381 -17467 -3347
rect -17433 -3381 -17420 -3347
rect -17480 -3419 -17420 -3381
rect -17480 -3453 -17467 -3419
rect -17433 -3453 -17420 -3419
rect -17480 -3491 -17420 -3453
rect -17480 -3525 -17467 -3491
rect -17433 -3525 -17420 -3491
rect -17480 -3563 -17420 -3525
rect -17480 -3597 -17467 -3563
rect -17433 -3597 -17420 -3563
rect -17480 -3635 -17420 -3597
rect -17480 -3669 -17467 -3635
rect -17433 -3669 -17420 -3635
rect -17480 -3707 -17420 -3669
rect -17480 -3741 -17467 -3707
rect -17433 -3741 -17420 -3707
rect -17480 -3779 -17420 -3741
rect -17480 -3813 -17467 -3779
rect -17433 -3813 -17420 -3779
rect -17480 -3851 -17420 -3813
rect -17480 -3885 -17467 -3851
rect -17433 -3885 -17420 -3851
rect -17480 -3923 -17420 -3885
rect -17480 -3957 -17467 -3923
rect -17433 -3957 -17420 -3923
rect -17480 -3995 -17420 -3957
rect -17480 -4029 -17467 -3995
rect -17433 -4029 -17420 -3995
rect -17480 -4067 -17420 -4029
rect -17480 -4101 -17467 -4067
rect -17433 -4101 -17420 -4067
rect -17480 -4139 -17420 -4101
rect -17480 -4173 -17467 -4139
rect -17433 -4173 -17420 -4139
rect -17480 -4211 -17420 -4173
rect -17480 -4245 -17467 -4211
rect -17433 -4245 -17420 -4211
rect -17480 -4283 -17420 -4245
rect -17480 -4317 -17467 -4283
rect -17433 -4317 -17420 -4283
rect -17480 -4355 -17420 -4317
rect -17480 -4380 -17467 -4355
rect -17500 -4389 -17467 -4380
rect -17433 -4380 -17420 -4355
rect 35320 -2771 35380 -2760
rect 35320 -2805 35333 -2771
rect 35367 -2805 35380 -2771
rect 35320 -2843 35380 -2805
rect 35320 -2877 35333 -2843
rect 35367 -2877 35380 -2843
rect 35320 -2915 35380 -2877
rect 35320 -2949 35333 -2915
rect 35367 -2949 35380 -2915
rect 35320 -2987 35380 -2949
rect 35320 -3021 35333 -2987
rect 35367 -3021 35380 -2987
rect 35320 -3059 35380 -3021
rect 35320 -3093 35333 -3059
rect 35367 -3093 35380 -3059
rect 35320 -3131 35380 -3093
rect 35320 -3165 35333 -3131
rect 35367 -3165 35380 -3131
rect 35320 -3203 35380 -3165
rect 35320 -3237 35333 -3203
rect 35367 -3237 35380 -3203
rect 35320 -3275 35380 -3237
rect 35320 -3309 35333 -3275
rect 35367 -3309 35380 -3275
rect 35320 -3347 35380 -3309
rect 35320 -3381 35333 -3347
rect 35367 -3381 35380 -3347
rect 35320 -3419 35380 -3381
rect 35320 -3453 35333 -3419
rect 35367 -3453 35380 -3419
rect 35320 -3491 35380 -3453
rect 35320 -3525 35333 -3491
rect 35367 -3525 35380 -3491
rect 35320 -3563 35380 -3525
rect 35320 -3597 35333 -3563
rect 35367 -3597 35380 -3563
rect 35320 -3635 35380 -3597
rect 35320 -3669 35333 -3635
rect 35367 -3669 35380 -3635
rect 35320 -3707 35380 -3669
rect 35320 -3741 35333 -3707
rect 35367 -3741 35380 -3707
rect 35320 -3779 35380 -3741
rect 35320 -3813 35333 -3779
rect 35367 -3813 35380 -3779
rect 35320 -3851 35380 -3813
rect 35320 -3885 35333 -3851
rect 35367 -3885 35380 -3851
rect 35320 -3923 35380 -3885
rect 35320 -3957 35333 -3923
rect 35367 -3957 35380 -3923
rect 35320 -3995 35380 -3957
rect 35320 -4029 35333 -3995
rect 35367 -4029 35380 -3995
rect 35320 -4067 35380 -4029
rect 35320 -4101 35333 -4067
rect 35367 -4101 35380 -4067
rect 35320 -4139 35380 -4101
rect 35320 -4173 35333 -4139
rect 35367 -4173 35380 -4139
rect 35320 -4211 35380 -4173
rect 35320 -4245 35333 -4211
rect 35367 -4245 35380 -4211
rect 35320 -4283 35380 -4245
rect 35320 -4317 35333 -4283
rect 35367 -4317 35380 -4283
rect 35320 -4355 35380 -4317
rect 35320 -4380 35333 -4355
rect -17433 -4389 35333 -4380
rect 35367 -4380 35380 -4355
rect 35367 -4389 35400 -4380
rect -17500 -4427 35400 -4389
rect -17500 -4440 -17467 -4427
rect -17480 -4461 -17467 -4440
rect -17433 -4440 35333 -4427
rect -17433 -4461 -17420 -4440
rect -17480 -4499 -17420 -4461
rect -17480 -4533 -17467 -4499
rect -17433 -4533 -17420 -4499
rect -17480 -4571 -17420 -4533
rect -17480 -4605 -17467 -4571
rect -17433 -4605 -17420 -4571
rect -17480 -4643 -17420 -4605
rect -17480 -4677 -17467 -4643
rect -17433 -4677 -17420 -4643
rect -17480 -4715 -17420 -4677
rect -17480 -4749 -17467 -4715
rect -17433 -4749 -17420 -4715
rect -17480 -4787 -17420 -4749
rect -17480 -4821 -17467 -4787
rect -17433 -4821 -17420 -4787
rect -17480 -4859 -17420 -4821
rect -17480 -4893 -17467 -4859
rect -17433 -4893 -17420 -4859
rect -17480 -4931 -17420 -4893
rect -17480 -4965 -17467 -4931
rect -17433 -4965 -17420 -4931
rect -17480 -5003 -17420 -4965
rect -17480 -5037 -17467 -5003
rect -17433 -5037 -17420 -5003
rect -17480 -5075 -17420 -5037
rect -17480 -5109 -17467 -5075
rect -17433 -5109 -17420 -5075
rect -17480 -5147 -17420 -5109
rect -17480 -5181 -17467 -5147
rect -17433 -5181 -17420 -5147
rect -17480 -5219 -17420 -5181
rect -17480 -5253 -17467 -5219
rect -17433 -5253 -17420 -5219
rect -17480 -5291 -17420 -5253
rect -17480 -5325 -17467 -5291
rect -17433 -5325 -17420 -5291
rect -17480 -5363 -17420 -5325
rect -17480 -5397 -17467 -5363
rect -17433 -5397 -17420 -5363
rect -17480 -5435 -17420 -5397
rect -17480 -5469 -17467 -5435
rect -17433 -5469 -17420 -5435
rect -17480 -5507 -17420 -5469
rect -17480 -5541 -17467 -5507
rect -17433 -5541 -17420 -5507
rect -17480 -5579 -17420 -5541
rect -17480 -5613 -17467 -5579
rect -17433 -5613 -17420 -5579
rect -17480 -5651 -17420 -5613
rect -17480 -5685 -17467 -5651
rect -17433 -5685 -17420 -5651
rect -17480 -5723 -17420 -5685
rect -17480 -5757 -17467 -5723
rect -17433 -5757 -17420 -5723
rect -17480 -5795 -17420 -5757
rect -17480 -5829 -17467 -5795
rect -17433 -5829 -17420 -5795
rect -17480 -5867 -17420 -5829
rect -17480 -5901 -17467 -5867
rect -17433 -5901 -17420 -5867
rect -17480 -5939 -17420 -5901
rect -17480 -5973 -17467 -5939
rect -17433 -5973 -17420 -5939
rect -17480 -6011 -17420 -5973
rect -17480 -6045 -17467 -6011
rect -17433 -6045 -17420 -6011
rect -17480 -6083 -17420 -6045
rect -17480 -6117 -17467 -6083
rect -17433 -6117 -17420 -6083
rect -17480 -6155 -17420 -6117
rect -17480 -6189 -17467 -6155
rect -17433 -6189 -17420 -6155
rect -17480 -6200 -17420 -6189
rect 35320 -4461 35333 -4440
rect 35367 -4440 35400 -4427
rect 35367 -4461 35380 -4440
rect 35320 -4499 35380 -4461
rect 35320 -4533 35333 -4499
rect 35367 -4533 35380 -4499
rect 35320 -4571 35380 -4533
rect 35320 -4605 35333 -4571
rect 35367 -4605 35380 -4571
rect 35320 -4643 35380 -4605
rect 35320 -4677 35333 -4643
rect 35367 -4677 35380 -4643
rect 35320 -4715 35380 -4677
rect 35320 -4749 35333 -4715
rect 35367 -4749 35380 -4715
rect 35320 -4787 35380 -4749
rect 35320 -4821 35333 -4787
rect 35367 -4821 35380 -4787
rect 35320 -4859 35380 -4821
rect 35320 -4893 35333 -4859
rect 35367 -4893 35380 -4859
rect 35320 -4931 35380 -4893
rect 35320 -4965 35333 -4931
rect 35367 -4965 35380 -4931
rect 35320 -5003 35380 -4965
rect 35320 -5037 35333 -5003
rect 35367 -5037 35380 -5003
rect 35320 -5075 35380 -5037
rect 35320 -5109 35333 -5075
rect 35367 -5109 35380 -5075
rect 35320 -5147 35380 -5109
rect 35320 -5181 35333 -5147
rect 35367 -5181 35380 -5147
rect 35320 -5219 35380 -5181
rect 35320 -5253 35333 -5219
rect 35367 -5253 35380 -5219
rect 35320 -5291 35380 -5253
rect 35320 -5325 35333 -5291
rect 35367 -5325 35380 -5291
rect 35320 -5363 35380 -5325
rect 35320 -5397 35333 -5363
rect 35367 -5397 35380 -5363
rect 35320 -5435 35380 -5397
rect 35320 -5469 35333 -5435
rect 35367 -5469 35380 -5435
rect 35320 -5507 35380 -5469
rect 35320 -5541 35333 -5507
rect 35367 -5541 35380 -5507
rect 35320 -5579 35380 -5541
rect 35320 -5613 35333 -5579
rect 35367 -5613 35380 -5579
rect 35320 -5651 35380 -5613
rect 35320 -5685 35333 -5651
rect 35367 -5685 35380 -5651
rect 35320 -5723 35380 -5685
rect 35320 -5757 35333 -5723
rect 35367 -5757 35380 -5723
rect 35320 -5795 35380 -5757
rect 35320 -5829 35333 -5795
rect 35367 -5829 35380 -5795
rect 35320 -5867 35380 -5829
rect 35320 -5901 35333 -5867
rect 35367 -5901 35380 -5867
rect 35320 -5939 35380 -5901
rect 35320 -5973 35333 -5939
rect 35367 -5973 35380 -5939
rect 35320 -6011 35380 -5973
rect 35320 -6045 35333 -6011
rect 35367 -6045 35380 -6011
rect 35320 -6083 35380 -6045
rect 35320 -6117 35333 -6083
rect 35367 -6117 35380 -6083
rect 35320 -6155 35380 -6117
rect 35320 -6189 35333 -6155
rect 35367 -6189 35380 -6155
rect 35320 -6200 35380 -6189
rect -17500 -6227 35400 -6200
rect -17500 -6260 -17467 -6227
rect -17480 -6261 -17467 -6260
rect -17433 -6260 35333 -6227
rect -17433 -6261 -17420 -6260
rect -17480 -6299 -17420 -6261
rect -17480 -6333 -17467 -6299
rect -17433 -6333 -17420 -6299
rect -17480 -6371 -17420 -6333
rect -17480 -6405 -17467 -6371
rect -17433 -6405 -17420 -6371
rect -17480 -6443 -17420 -6405
rect -17480 -6477 -17467 -6443
rect -17433 -6477 -17420 -6443
rect -17480 -6515 -17420 -6477
rect -17480 -6549 -17467 -6515
rect -17433 -6549 -17420 -6515
rect -17480 -6587 -17420 -6549
rect -17480 -6621 -17467 -6587
rect -17433 -6621 -17420 -6587
rect -17480 -6659 -17420 -6621
rect -17480 -6693 -17467 -6659
rect -17433 -6693 -17420 -6659
rect -17480 -6731 -17420 -6693
rect -17480 -6765 -17467 -6731
rect -17433 -6765 -17420 -6731
rect -17480 -6803 -17420 -6765
rect -17480 -6837 -17467 -6803
rect -17433 -6837 -17420 -6803
rect -17480 -6875 -17420 -6837
rect -17480 -6909 -17467 -6875
rect -17433 -6909 -17420 -6875
rect -17480 -6947 -17420 -6909
rect -17480 -6981 -17467 -6947
rect -17433 -6981 -17420 -6947
rect -17480 -7019 -17420 -6981
rect -17480 -7053 -17467 -7019
rect -17433 -7053 -17420 -7019
rect -17480 -7091 -17420 -7053
rect -17480 -7125 -17467 -7091
rect -17433 -7125 -17420 -7091
rect -17480 -7163 -17420 -7125
rect -17480 -7197 -17467 -7163
rect -17433 -7197 -17420 -7163
rect -17480 -7200 -17420 -7197
rect 35320 -6261 35333 -6260
rect 35367 -6260 35400 -6227
rect 35367 -6261 35380 -6260
rect 35320 -6299 35380 -6261
rect 35320 -6333 35333 -6299
rect 35367 -6333 35380 -6299
rect 35320 -6371 35380 -6333
rect 35320 -6405 35333 -6371
rect 35367 -6405 35380 -6371
rect 35320 -6443 35380 -6405
rect 35320 -6477 35333 -6443
rect 35367 -6477 35380 -6443
rect 35320 -6515 35380 -6477
rect 35320 -6549 35333 -6515
rect 35367 -6549 35380 -6515
rect 35320 -6587 35380 -6549
rect 35320 -6621 35333 -6587
rect 35367 -6621 35380 -6587
rect 35320 -6659 35380 -6621
rect 35320 -6693 35333 -6659
rect 35367 -6693 35380 -6659
rect 35320 -6731 35380 -6693
rect 35320 -6765 35333 -6731
rect 35367 -6765 35380 -6731
rect 35320 -6803 35380 -6765
rect 35320 -6837 35333 -6803
rect 35367 -6837 35380 -6803
rect 35320 -6875 35380 -6837
rect 35320 -6909 35333 -6875
rect 35367 -6909 35380 -6875
rect 35320 -6947 35380 -6909
rect 35320 -6981 35333 -6947
rect 35367 -6981 35380 -6947
rect 35320 -7019 35380 -6981
rect 35320 -7053 35333 -7019
rect 35367 -7053 35380 -7019
rect 35320 -7091 35380 -7053
rect 35320 -7125 35333 -7091
rect 35367 -7125 35380 -7091
rect 35320 -7163 35380 -7125
rect 35320 -7197 35333 -7163
rect 35367 -7197 35380 -7163
rect 35320 -7200 35380 -7197
rect -17340 -7233 35220 -7220
rect -17340 -7267 -17321 -7233
rect -17287 -7267 -17249 -7233
rect -17215 -7267 -17177 -7233
rect -17143 -7267 -17105 -7233
rect -17071 -7267 -17033 -7233
rect -16999 -7267 -16961 -7233
rect -16927 -7267 -16889 -7233
rect -16855 -7267 -16817 -7233
rect -16783 -7267 -16745 -7233
rect -16711 -7267 -16673 -7233
rect -16639 -7267 -16601 -7233
rect -16567 -7267 -16529 -7233
rect -16495 -7267 -16457 -7233
rect -16423 -7267 -16385 -7233
rect -16351 -7267 -16313 -7233
rect -16279 -7267 -16241 -7233
rect -16207 -7267 -16169 -7233
rect -16135 -7267 -16097 -7233
rect -16063 -7267 -16025 -7233
rect -15991 -7267 -15953 -7233
rect -15919 -7267 -15881 -7233
rect -15847 -7267 -15809 -7233
rect -15775 -7267 -15737 -7233
rect -15703 -7267 -15665 -7233
rect -15631 -7267 -15593 -7233
rect -15559 -7267 -15521 -7233
rect -15487 -7267 -15449 -7233
rect -15415 -7267 -15377 -7233
rect -15343 -7267 -15305 -7233
rect -15271 -7267 -15233 -7233
rect -15199 -7267 -15161 -7233
rect -15127 -7267 -15089 -7233
rect -15055 -7267 -15017 -7233
rect -14983 -7267 -14945 -7233
rect -14911 -7267 -14873 -7233
rect -14839 -7267 -14801 -7233
rect -14767 -7267 -14729 -7233
rect -14695 -7267 -14657 -7233
rect -14623 -7267 -14585 -7233
rect -14551 -7267 -14513 -7233
rect -14479 -7267 -14441 -7233
rect -14407 -7267 -14369 -7233
rect -14335 -7267 -14297 -7233
rect -14263 -7267 -14225 -7233
rect -14191 -7267 -14153 -7233
rect -14119 -7267 -14081 -7233
rect -14047 -7267 -14009 -7233
rect -13975 -7267 -13937 -7233
rect -13903 -7267 -13865 -7233
rect -13831 -7267 -13793 -7233
rect -13759 -7267 -13721 -7233
rect -13687 -7267 -13649 -7233
rect -13615 -7267 -13577 -7233
rect -13543 -7267 -13505 -7233
rect -13471 -7267 -13433 -7233
rect -13399 -7267 -13361 -7233
rect -13327 -7267 -13289 -7233
rect -13255 -7267 -13217 -7233
rect -13183 -7267 -13145 -7233
rect -13111 -7267 -13073 -7233
rect -13039 -7267 -13001 -7233
rect -12967 -7267 -12929 -7233
rect -12895 -7267 -12857 -7233
rect -12823 -7267 -12785 -7233
rect -12751 -7267 -12713 -7233
rect -12679 -7267 -12641 -7233
rect -12607 -7267 -12569 -7233
rect -12535 -7267 -12497 -7233
rect -12463 -7267 -12425 -7233
rect -12391 -7267 -12353 -7233
rect -12319 -7267 -12281 -7233
rect -12247 -7267 -12209 -7233
rect -12175 -7267 -12137 -7233
rect -12103 -7267 -12065 -7233
rect -12031 -7267 -11993 -7233
rect -11959 -7267 -11921 -7233
rect -11887 -7267 -11849 -7233
rect -11815 -7267 -11777 -7233
rect -11743 -7267 -11705 -7233
rect -11671 -7267 -11633 -7233
rect -11599 -7267 -11561 -7233
rect -11527 -7267 -11489 -7233
rect -11455 -7267 -11417 -7233
rect -11383 -7267 -11345 -7233
rect -11311 -7267 -11273 -7233
rect -11239 -7267 -11201 -7233
rect -11167 -7267 -11129 -7233
rect -11095 -7267 -11057 -7233
rect -11023 -7267 -10985 -7233
rect -10951 -7267 -10913 -7233
rect -10879 -7267 -10841 -7233
rect -10807 -7267 -10769 -7233
rect -10735 -7267 -10697 -7233
rect -10663 -7267 -10625 -7233
rect -10591 -7267 -10553 -7233
rect -10519 -7267 -10481 -7233
rect -10447 -7267 -10409 -7233
rect -10375 -7267 -10337 -7233
rect -10303 -7267 -10265 -7233
rect -10231 -7267 -10193 -7233
rect -10159 -7267 -10121 -7233
rect -10087 -7267 -10049 -7233
rect -10015 -7267 -9977 -7233
rect -9943 -7267 -9905 -7233
rect -9871 -7267 -9833 -7233
rect -9799 -7267 -9761 -7233
rect -9727 -7267 -9689 -7233
rect -9655 -7267 -9617 -7233
rect -9583 -7267 -9545 -7233
rect -9511 -7267 -9473 -7233
rect -9439 -7267 -9401 -7233
rect -9367 -7267 -9329 -7233
rect -9295 -7267 -9257 -7233
rect -9223 -7267 -9185 -7233
rect -9151 -7267 -9113 -7233
rect -9079 -7267 -9041 -7233
rect -9007 -7267 -8969 -7233
rect -8935 -7267 -8897 -7233
rect -8863 -7267 -8825 -7233
rect -8791 -7267 -8753 -7233
rect -8719 -7267 -8681 -7233
rect -8647 -7267 -8609 -7233
rect -8575 -7267 -8537 -7233
rect -8503 -7267 -8465 -7233
rect -8431 -7267 -8393 -7233
rect -8359 -7267 -8321 -7233
rect -8287 -7267 -8249 -7233
rect -8215 -7267 -8177 -7233
rect -8143 -7267 -8105 -7233
rect -8071 -7267 -8033 -7233
rect -7999 -7267 -7961 -7233
rect -7927 -7267 -7889 -7233
rect -7855 -7267 -7817 -7233
rect -7783 -7267 -7745 -7233
rect -7711 -7267 -7673 -7233
rect -7639 -7267 -7601 -7233
rect -7567 -7267 -7529 -7233
rect -7495 -7267 -7457 -7233
rect -7423 -7267 -7385 -7233
rect -7351 -7267 -7313 -7233
rect -7279 -7267 -7241 -7233
rect -7207 -7267 -7169 -7233
rect -7135 -7267 -7097 -7233
rect -7063 -7267 -7025 -7233
rect -6991 -7267 -6953 -7233
rect -6919 -7267 -6881 -7233
rect -6847 -7267 -6809 -7233
rect -6775 -7267 -6737 -7233
rect -6703 -7267 -6665 -7233
rect -6631 -7267 -6593 -7233
rect -6559 -7267 -6521 -7233
rect -6487 -7267 -6449 -7233
rect -6415 -7267 -6377 -7233
rect -6343 -7267 -6305 -7233
rect -6271 -7267 -6233 -7233
rect -6199 -7267 -6161 -7233
rect -6127 -7267 -6089 -7233
rect -6055 -7267 -6017 -7233
rect -5983 -7267 -5945 -7233
rect -5911 -7267 -5873 -7233
rect -5839 -7267 -5801 -7233
rect -5767 -7267 -5729 -7233
rect -5695 -7267 -5657 -7233
rect -5623 -7267 -5585 -7233
rect -5551 -7267 -5513 -7233
rect -5479 -7267 -5441 -7233
rect -5407 -7267 -5369 -7233
rect -5335 -7267 -5297 -7233
rect -5263 -7267 -5225 -7233
rect -5191 -7267 -5153 -7233
rect -5119 -7267 -5081 -7233
rect -5047 -7267 -5009 -7233
rect -4975 -7267 -4937 -7233
rect -4903 -7267 -4865 -7233
rect -4831 -7267 -4793 -7233
rect -4759 -7267 -4721 -7233
rect -4687 -7267 -4649 -7233
rect -4615 -7267 -4577 -7233
rect -4543 -7267 -4505 -7233
rect -4471 -7267 -4433 -7233
rect -4399 -7267 -4361 -7233
rect -4327 -7267 -4289 -7233
rect -4255 -7267 -4217 -7233
rect -4183 -7267 -4145 -7233
rect -4111 -7267 -4073 -7233
rect -4039 -7267 -4001 -7233
rect -3967 -7267 -3929 -7233
rect -3895 -7267 -3857 -7233
rect -3823 -7267 -3785 -7233
rect -3751 -7267 -3713 -7233
rect -3679 -7267 -3641 -7233
rect -3607 -7267 -3569 -7233
rect -3535 -7267 -3497 -7233
rect -3463 -7267 -3425 -7233
rect -3391 -7267 -3353 -7233
rect -3319 -7267 -3281 -7233
rect -3247 -7267 -3209 -7233
rect -3175 -7267 -3137 -7233
rect -3103 -7267 -3065 -7233
rect -3031 -7267 -2993 -7233
rect -2959 -7267 -2921 -7233
rect -2887 -7267 -2849 -7233
rect -2815 -7267 -2777 -7233
rect -2743 -7267 -2705 -7233
rect -2671 -7267 -2633 -7233
rect -2599 -7267 -2561 -7233
rect -2527 -7267 -2489 -7233
rect -2455 -7267 -2417 -7233
rect -2383 -7267 -2345 -7233
rect -2311 -7267 -2273 -7233
rect -2239 -7267 -2201 -7233
rect -2167 -7267 -2129 -7233
rect -2095 -7267 -2057 -7233
rect -2023 -7267 -1985 -7233
rect -1951 -7267 -1913 -7233
rect -1879 -7267 -1841 -7233
rect -1807 -7267 -1769 -7233
rect -1735 -7267 -1697 -7233
rect -1663 -7267 -1625 -7233
rect -1591 -7267 -1553 -7233
rect -1519 -7267 -1481 -7233
rect -1447 -7267 -1409 -7233
rect -1375 -7267 -1337 -7233
rect -1303 -7267 -1265 -7233
rect -1231 -7267 -1193 -7233
rect -1159 -7267 -1121 -7233
rect -1087 -7267 -1049 -7233
rect -1015 -7267 -977 -7233
rect -943 -7267 -905 -7233
rect -871 -7267 -833 -7233
rect -799 -7267 -761 -7233
rect -727 -7267 -689 -7233
rect -655 -7267 -617 -7233
rect -583 -7267 -545 -7233
rect -511 -7267 -473 -7233
rect -439 -7267 -401 -7233
rect -367 -7267 -329 -7233
rect -295 -7267 -257 -7233
rect -223 -7267 -185 -7233
rect -151 -7267 -113 -7233
rect -79 -7267 -41 -7233
rect -7 -7267 31 -7233
rect 65 -7267 103 -7233
rect 137 -7267 175 -7233
rect 209 -7267 247 -7233
rect 281 -7267 319 -7233
rect 353 -7267 391 -7233
rect 425 -7267 463 -7233
rect 497 -7267 535 -7233
rect 569 -7267 607 -7233
rect 641 -7267 679 -7233
rect 713 -7267 751 -7233
rect 785 -7267 823 -7233
rect 857 -7267 895 -7233
rect 929 -7267 967 -7233
rect 1001 -7267 1039 -7233
rect 1073 -7267 1111 -7233
rect 1145 -7267 1183 -7233
rect 1217 -7267 1255 -7233
rect 1289 -7267 1327 -7233
rect 1361 -7267 1399 -7233
rect 1433 -7267 1471 -7233
rect 1505 -7267 1543 -7233
rect 1577 -7267 1615 -7233
rect 1649 -7267 1687 -7233
rect 1721 -7267 1759 -7233
rect 1793 -7267 1831 -7233
rect 1865 -7267 1903 -7233
rect 1937 -7267 1975 -7233
rect 2009 -7267 2047 -7233
rect 2081 -7267 2119 -7233
rect 2153 -7267 2191 -7233
rect 2225 -7267 2263 -7233
rect 2297 -7267 2335 -7233
rect 2369 -7267 2407 -7233
rect 2441 -7267 2479 -7233
rect 2513 -7267 2551 -7233
rect 2585 -7267 2623 -7233
rect 2657 -7267 2695 -7233
rect 2729 -7267 2767 -7233
rect 2801 -7267 2839 -7233
rect 2873 -7267 2911 -7233
rect 2945 -7267 2983 -7233
rect 3017 -7267 3055 -7233
rect 3089 -7267 3127 -7233
rect 3161 -7267 3199 -7233
rect 3233 -7267 3271 -7233
rect 3305 -7267 3343 -7233
rect 3377 -7267 3415 -7233
rect 3449 -7267 3487 -7233
rect 3521 -7267 3559 -7233
rect 3593 -7267 3631 -7233
rect 3665 -7267 3703 -7233
rect 3737 -7267 3775 -7233
rect 3809 -7267 3847 -7233
rect 3881 -7267 3919 -7233
rect 3953 -7267 3991 -7233
rect 4025 -7267 4063 -7233
rect 4097 -7267 4135 -7233
rect 4169 -7267 4207 -7233
rect 4241 -7267 4279 -7233
rect 4313 -7267 4351 -7233
rect 4385 -7267 4423 -7233
rect 4457 -7267 4495 -7233
rect 4529 -7267 4567 -7233
rect 4601 -7267 4639 -7233
rect 4673 -7267 4711 -7233
rect 4745 -7267 4783 -7233
rect 4817 -7267 4855 -7233
rect 4889 -7267 4927 -7233
rect 4961 -7267 4999 -7233
rect 5033 -7267 5071 -7233
rect 5105 -7267 5143 -7233
rect 5177 -7267 5215 -7233
rect 5249 -7267 5287 -7233
rect 5321 -7267 5359 -7233
rect 5393 -7267 5431 -7233
rect 5465 -7267 5503 -7233
rect 5537 -7267 5575 -7233
rect 5609 -7267 5647 -7233
rect 5681 -7267 5719 -7233
rect 5753 -7267 5791 -7233
rect 5825 -7267 5863 -7233
rect 5897 -7267 5935 -7233
rect 5969 -7267 6007 -7233
rect 6041 -7267 6079 -7233
rect 6113 -7267 6151 -7233
rect 6185 -7267 6223 -7233
rect 6257 -7267 6295 -7233
rect 6329 -7267 6367 -7233
rect 6401 -7267 6439 -7233
rect 6473 -7267 6511 -7233
rect 6545 -7267 6583 -7233
rect 6617 -7267 6655 -7233
rect 6689 -7267 6727 -7233
rect 6761 -7267 6799 -7233
rect 6833 -7267 6871 -7233
rect 6905 -7267 6943 -7233
rect 6977 -7267 7015 -7233
rect 7049 -7267 7087 -7233
rect 7121 -7267 7159 -7233
rect 7193 -7267 7231 -7233
rect 7265 -7267 7303 -7233
rect 7337 -7267 7375 -7233
rect 7409 -7267 7447 -7233
rect 7481 -7267 7519 -7233
rect 7553 -7267 7591 -7233
rect 7625 -7267 7663 -7233
rect 7697 -7267 7735 -7233
rect 7769 -7267 7807 -7233
rect 7841 -7267 7879 -7233
rect 7913 -7267 7951 -7233
rect 7985 -7267 8023 -7233
rect 8057 -7267 8095 -7233
rect 8129 -7267 8167 -7233
rect 8201 -7267 8239 -7233
rect 8273 -7267 8311 -7233
rect 8345 -7267 8383 -7233
rect 8417 -7267 8455 -7233
rect 8489 -7267 8527 -7233
rect 8561 -7267 8599 -7233
rect 8633 -7267 8671 -7233
rect 8705 -7267 8743 -7233
rect 8777 -7267 8815 -7233
rect 8849 -7267 8887 -7233
rect 8921 -7267 8959 -7233
rect 8993 -7267 9031 -7233
rect 9065 -7267 9103 -7233
rect 9137 -7267 9175 -7233
rect 9209 -7267 9247 -7233
rect 9281 -7267 9319 -7233
rect 9353 -7267 9391 -7233
rect 9425 -7267 9463 -7233
rect 9497 -7267 9535 -7233
rect 9569 -7267 9607 -7233
rect 9641 -7267 9679 -7233
rect 9713 -7267 9751 -7233
rect 9785 -7267 9823 -7233
rect 9857 -7267 9895 -7233
rect 9929 -7267 9967 -7233
rect 10001 -7267 10039 -7233
rect 10073 -7267 10111 -7233
rect 10145 -7267 10183 -7233
rect 10217 -7267 10255 -7233
rect 10289 -7267 10327 -7233
rect 10361 -7267 10399 -7233
rect 10433 -7267 10471 -7233
rect 10505 -7267 10543 -7233
rect 10577 -7267 10615 -7233
rect 10649 -7267 10687 -7233
rect 10721 -7267 10759 -7233
rect 10793 -7267 10831 -7233
rect 10865 -7267 10903 -7233
rect 10937 -7267 10975 -7233
rect 11009 -7267 11047 -7233
rect 11081 -7267 11119 -7233
rect 11153 -7267 11191 -7233
rect 11225 -7267 11263 -7233
rect 11297 -7267 11335 -7233
rect 11369 -7267 11407 -7233
rect 11441 -7267 11479 -7233
rect 11513 -7267 11551 -7233
rect 11585 -7267 11623 -7233
rect 11657 -7267 11695 -7233
rect 11729 -7267 11767 -7233
rect 11801 -7267 11839 -7233
rect 11873 -7267 11911 -7233
rect 11945 -7267 11983 -7233
rect 12017 -7267 12055 -7233
rect 12089 -7267 12127 -7233
rect 12161 -7267 12199 -7233
rect 12233 -7267 12271 -7233
rect 12305 -7267 12343 -7233
rect 12377 -7267 12415 -7233
rect 12449 -7267 12487 -7233
rect 12521 -7267 12559 -7233
rect 12593 -7267 12631 -7233
rect 12665 -7267 12703 -7233
rect 12737 -7267 12775 -7233
rect 12809 -7267 12847 -7233
rect 12881 -7267 12919 -7233
rect 12953 -7267 12991 -7233
rect 13025 -7267 13063 -7233
rect 13097 -7267 13135 -7233
rect 13169 -7267 13207 -7233
rect 13241 -7267 13279 -7233
rect 13313 -7267 13351 -7233
rect 13385 -7267 13423 -7233
rect 13457 -7267 13495 -7233
rect 13529 -7267 13567 -7233
rect 13601 -7267 13639 -7233
rect 13673 -7267 13711 -7233
rect 13745 -7267 13783 -7233
rect 13817 -7267 13855 -7233
rect 13889 -7267 13927 -7233
rect 13961 -7267 13999 -7233
rect 14033 -7267 14071 -7233
rect 14105 -7267 14143 -7233
rect 14177 -7267 14215 -7233
rect 14249 -7267 14287 -7233
rect 14321 -7267 14359 -7233
rect 14393 -7267 14431 -7233
rect 14465 -7267 14503 -7233
rect 14537 -7267 14575 -7233
rect 14609 -7267 14647 -7233
rect 14681 -7267 14719 -7233
rect 14753 -7267 14791 -7233
rect 14825 -7267 14863 -7233
rect 14897 -7267 14935 -7233
rect 14969 -7267 15007 -7233
rect 15041 -7267 15079 -7233
rect 15113 -7267 15151 -7233
rect 15185 -7267 15223 -7233
rect 15257 -7267 15295 -7233
rect 15329 -7267 15367 -7233
rect 15401 -7267 15439 -7233
rect 15473 -7267 15511 -7233
rect 15545 -7267 15583 -7233
rect 15617 -7267 15655 -7233
rect 15689 -7267 15727 -7233
rect 15761 -7267 15799 -7233
rect 15833 -7267 15871 -7233
rect 15905 -7267 15943 -7233
rect 15977 -7267 16015 -7233
rect 16049 -7267 16087 -7233
rect 16121 -7267 16159 -7233
rect 16193 -7267 16231 -7233
rect 16265 -7267 16303 -7233
rect 16337 -7267 16375 -7233
rect 16409 -7267 16447 -7233
rect 16481 -7267 16519 -7233
rect 16553 -7267 16591 -7233
rect 16625 -7267 16663 -7233
rect 16697 -7267 16735 -7233
rect 16769 -7267 16807 -7233
rect 16841 -7267 16879 -7233
rect 16913 -7267 16951 -7233
rect 16985 -7267 17023 -7233
rect 17057 -7267 17095 -7233
rect 17129 -7267 17167 -7233
rect 17201 -7267 17239 -7233
rect 17273 -7267 17311 -7233
rect 17345 -7267 17383 -7233
rect 17417 -7267 17455 -7233
rect 17489 -7267 17527 -7233
rect 17561 -7267 17599 -7233
rect 17633 -7267 17671 -7233
rect 17705 -7267 17743 -7233
rect 17777 -7267 17815 -7233
rect 17849 -7267 17887 -7233
rect 17921 -7267 17959 -7233
rect 17993 -7267 18031 -7233
rect 18065 -7267 18103 -7233
rect 18137 -7267 18175 -7233
rect 18209 -7267 18247 -7233
rect 18281 -7267 18319 -7233
rect 18353 -7267 18391 -7233
rect 18425 -7267 18463 -7233
rect 18497 -7267 18535 -7233
rect 18569 -7267 18607 -7233
rect 18641 -7267 18679 -7233
rect 18713 -7267 18751 -7233
rect 18785 -7267 18823 -7233
rect 18857 -7267 18895 -7233
rect 18929 -7267 18967 -7233
rect 19001 -7267 19039 -7233
rect 19073 -7267 19111 -7233
rect 19145 -7267 19183 -7233
rect 19217 -7267 19255 -7233
rect 19289 -7267 19327 -7233
rect 19361 -7267 19399 -7233
rect 19433 -7267 19471 -7233
rect 19505 -7267 19543 -7233
rect 19577 -7267 19615 -7233
rect 19649 -7267 19687 -7233
rect 19721 -7267 19759 -7233
rect 19793 -7267 19831 -7233
rect 19865 -7267 19903 -7233
rect 19937 -7267 19975 -7233
rect 20009 -7267 20047 -7233
rect 20081 -7267 20119 -7233
rect 20153 -7267 20191 -7233
rect 20225 -7267 20263 -7233
rect 20297 -7267 20335 -7233
rect 20369 -7267 20407 -7233
rect 20441 -7267 20479 -7233
rect 20513 -7267 20551 -7233
rect 20585 -7267 20623 -7233
rect 20657 -7267 20695 -7233
rect 20729 -7267 20767 -7233
rect 20801 -7267 20839 -7233
rect 20873 -7267 20911 -7233
rect 20945 -7267 20983 -7233
rect 21017 -7267 21055 -7233
rect 21089 -7267 21127 -7233
rect 21161 -7267 21199 -7233
rect 21233 -7267 21271 -7233
rect 21305 -7267 21343 -7233
rect 21377 -7267 21415 -7233
rect 21449 -7267 21487 -7233
rect 21521 -7267 21559 -7233
rect 21593 -7267 21631 -7233
rect 21665 -7267 21703 -7233
rect 21737 -7267 21775 -7233
rect 21809 -7267 21847 -7233
rect 21881 -7267 21919 -7233
rect 21953 -7267 21991 -7233
rect 22025 -7267 22063 -7233
rect 22097 -7267 22135 -7233
rect 22169 -7267 22207 -7233
rect 22241 -7267 22279 -7233
rect 22313 -7267 22351 -7233
rect 22385 -7267 22423 -7233
rect 22457 -7267 22495 -7233
rect 22529 -7267 22567 -7233
rect 22601 -7267 22639 -7233
rect 22673 -7267 22711 -7233
rect 22745 -7267 22783 -7233
rect 22817 -7267 22855 -7233
rect 22889 -7267 22927 -7233
rect 22961 -7267 22999 -7233
rect 23033 -7267 23071 -7233
rect 23105 -7267 23143 -7233
rect 23177 -7267 23215 -7233
rect 23249 -7267 23287 -7233
rect 23321 -7267 23359 -7233
rect 23393 -7267 23431 -7233
rect 23465 -7267 23503 -7233
rect 23537 -7267 23575 -7233
rect 23609 -7267 23647 -7233
rect 23681 -7267 23719 -7233
rect 23753 -7267 23791 -7233
rect 23825 -7267 23863 -7233
rect 23897 -7267 23935 -7233
rect 23969 -7267 24007 -7233
rect 24041 -7267 24079 -7233
rect 24113 -7267 24151 -7233
rect 24185 -7267 24223 -7233
rect 24257 -7267 24295 -7233
rect 24329 -7267 24367 -7233
rect 24401 -7267 24439 -7233
rect 24473 -7267 24511 -7233
rect 24545 -7267 24583 -7233
rect 24617 -7267 24655 -7233
rect 24689 -7267 24727 -7233
rect 24761 -7267 24799 -7233
rect 24833 -7267 24871 -7233
rect 24905 -7267 24943 -7233
rect 24977 -7267 25015 -7233
rect 25049 -7267 25087 -7233
rect 25121 -7267 25159 -7233
rect 25193 -7267 25231 -7233
rect 25265 -7267 25303 -7233
rect 25337 -7267 25375 -7233
rect 25409 -7267 25447 -7233
rect 25481 -7267 25519 -7233
rect 25553 -7267 25591 -7233
rect 25625 -7267 25663 -7233
rect 25697 -7267 25735 -7233
rect 25769 -7267 25807 -7233
rect 25841 -7267 25879 -7233
rect 25913 -7267 25951 -7233
rect 25985 -7267 26023 -7233
rect 26057 -7267 26095 -7233
rect 26129 -7267 26167 -7233
rect 26201 -7267 26239 -7233
rect 26273 -7267 26311 -7233
rect 26345 -7267 26383 -7233
rect 26417 -7267 26455 -7233
rect 26489 -7267 26527 -7233
rect 26561 -7267 26599 -7233
rect 26633 -7267 26671 -7233
rect 26705 -7267 26743 -7233
rect 26777 -7267 26815 -7233
rect 26849 -7267 26887 -7233
rect 26921 -7267 26959 -7233
rect 26993 -7267 27031 -7233
rect 27065 -7267 27103 -7233
rect 27137 -7267 27175 -7233
rect 27209 -7267 27247 -7233
rect 27281 -7267 27319 -7233
rect 27353 -7267 27391 -7233
rect 27425 -7267 27463 -7233
rect 27497 -7267 27535 -7233
rect 27569 -7267 27607 -7233
rect 27641 -7267 27679 -7233
rect 27713 -7267 27751 -7233
rect 27785 -7267 27823 -7233
rect 27857 -7267 27895 -7233
rect 27929 -7267 27967 -7233
rect 28001 -7267 28039 -7233
rect 28073 -7267 28111 -7233
rect 28145 -7267 28183 -7233
rect 28217 -7267 28255 -7233
rect 28289 -7267 28327 -7233
rect 28361 -7267 28399 -7233
rect 28433 -7267 28471 -7233
rect 28505 -7267 28543 -7233
rect 28577 -7267 28615 -7233
rect 28649 -7267 28687 -7233
rect 28721 -7267 28759 -7233
rect 28793 -7267 28831 -7233
rect 28865 -7267 28903 -7233
rect 28937 -7267 28975 -7233
rect 29009 -7267 29047 -7233
rect 29081 -7267 29119 -7233
rect 29153 -7267 29191 -7233
rect 29225 -7267 29263 -7233
rect 29297 -7267 29335 -7233
rect 29369 -7267 29407 -7233
rect 29441 -7267 29479 -7233
rect 29513 -7267 29551 -7233
rect 29585 -7267 29623 -7233
rect 29657 -7267 29695 -7233
rect 29729 -7267 29767 -7233
rect 29801 -7267 29839 -7233
rect 29873 -7267 29911 -7233
rect 29945 -7267 29983 -7233
rect 30017 -7267 30055 -7233
rect 30089 -7267 30127 -7233
rect 30161 -7267 30199 -7233
rect 30233 -7267 30271 -7233
rect 30305 -7267 30343 -7233
rect 30377 -7267 30415 -7233
rect 30449 -7267 30487 -7233
rect 30521 -7267 30559 -7233
rect 30593 -7267 30631 -7233
rect 30665 -7267 30703 -7233
rect 30737 -7267 30775 -7233
rect 30809 -7267 30847 -7233
rect 30881 -7267 30919 -7233
rect 30953 -7267 30991 -7233
rect 31025 -7267 31063 -7233
rect 31097 -7267 31135 -7233
rect 31169 -7267 31207 -7233
rect 31241 -7267 31279 -7233
rect 31313 -7267 31351 -7233
rect 31385 -7267 31423 -7233
rect 31457 -7267 31495 -7233
rect 31529 -7267 31567 -7233
rect 31601 -7267 31639 -7233
rect 31673 -7267 31711 -7233
rect 31745 -7267 31783 -7233
rect 31817 -7267 31855 -7233
rect 31889 -7267 31927 -7233
rect 31961 -7267 31999 -7233
rect 32033 -7267 32071 -7233
rect 32105 -7267 32143 -7233
rect 32177 -7267 32215 -7233
rect 32249 -7267 32287 -7233
rect 32321 -7267 32359 -7233
rect 32393 -7267 32431 -7233
rect 32465 -7267 32503 -7233
rect 32537 -7267 32575 -7233
rect 32609 -7267 32647 -7233
rect 32681 -7267 32719 -7233
rect 32753 -7267 32791 -7233
rect 32825 -7267 32863 -7233
rect 32897 -7267 32935 -7233
rect 32969 -7267 33007 -7233
rect 33041 -7267 33079 -7233
rect 33113 -7267 33151 -7233
rect 33185 -7267 33223 -7233
rect 33257 -7267 33295 -7233
rect 33329 -7267 33367 -7233
rect 33401 -7267 33439 -7233
rect 33473 -7267 33511 -7233
rect 33545 -7267 33583 -7233
rect 33617 -7267 33655 -7233
rect 33689 -7267 33727 -7233
rect 33761 -7267 33799 -7233
rect 33833 -7267 33871 -7233
rect 33905 -7267 33943 -7233
rect 33977 -7267 34015 -7233
rect 34049 -7267 34087 -7233
rect 34121 -7267 34159 -7233
rect 34193 -7267 34231 -7233
rect 34265 -7267 34303 -7233
rect 34337 -7267 34375 -7233
rect 34409 -7267 34447 -7233
rect 34481 -7267 34519 -7233
rect 34553 -7267 34591 -7233
rect 34625 -7267 34663 -7233
rect 34697 -7267 34735 -7233
rect 34769 -7267 34807 -7233
rect 34841 -7267 34879 -7233
rect 34913 -7267 34951 -7233
rect 34985 -7267 35023 -7233
rect 35057 -7267 35095 -7233
rect 35129 -7267 35167 -7233
rect 35201 -7267 35220 -7233
rect -17340 -7280 35220 -7267
<< viali >>
rect -17301 14833 -17267 14867
rect -17229 14833 -17195 14867
rect -17157 14833 -17123 14867
rect -17085 14833 -17051 14867
rect -17013 14833 -16979 14867
rect -16941 14833 -16907 14867
rect -16869 14833 -16835 14867
rect -16797 14833 -16763 14867
rect -16725 14833 -16691 14867
rect -16653 14833 -16619 14867
rect -16581 14833 -16547 14867
rect -16509 14833 -16475 14867
rect -16437 14833 -16403 14867
rect -16365 14833 -16331 14867
rect -16293 14833 -16259 14867
rect -16221 14833 -16187 14867
rect -16149 14833 -16115 14867
rect -16077 14833 -16043 14867
rect -16005 14833 -15971 14867
rect -15933 14833 -15899 14867
rect -15861 14833 -15827 14867
rect -15789 14833 -15755 14867
rect -15717 14833 -15683 14867
rect -15645 14833 -15611 14867
rect -15573 14833 -15539 14867
rect -15501 14833 -15467 14867
rect -15429 14833 -15395 14867
rect -15357 14833 -15323 14867
rect -15285 14833 -15251 14867
rect -15213 14833 -15179 14867
rect -15141 14833 -15107 14867
rect -15069 14833 -15035 14867
rect -14997 14833 -14963 14867
rect -14925 14833 -14891 14867
rect -14853 14833 -14819 14867
rect -14781 14833 -14747 14867
rect -14709 14833 -14675 14867
rect -14637 14833 -14603 14867
rect -14565 14833 -14531 14867
rect -14493 14833 -14459 14867
rect -14421 14833 -14387 14867
rect -14349 14833 -14315 14867
rect -14277 14833 -14243 14867
rect -14205 14833 -14171 14867
rect -14133 14833 -14099 14867
rect -14061 14833 -14027 14867
rect -13989 14833 -13955 14867
rect -13917 14833 -13883 14867
rect -13845 14833 -13811 14867
rect -13773 14833 -13739 14867
rect -13701 14833 -13667 14867
rect -13629 14833 -13595 14867
rect -13557 14833 -13523 14867
rect -13485 14833 -13451 14867
rect -13413 14833 -13379 14867
rect -13341 14833 -13307 14867
rect -13269 14833 -13235 14867
rect -13197 14833 -13163 14867
rect -13125 14833 -13091 14867
rect -13053 14833 -13019 14867
rect -12981 14833 -12947 14867
rect -12909 14833 -12875 14867
rect -12837 14833 -12803 14867
rect -12765 14833 -12731 14867
rect -12693 14833 -12659 14867
rect -12621 14833 -12587 14867
rect -12549 14833 -12515 14867
rect -12477 14833 -12443 14867
rect -12405 14833 -12371 14867
rect -12333 14833 -12299 14867
rect -12261 14833 -12227 14867
rect -12189 14833 -12155 14867
rect -12117 14833 -12083 14867
rect -12045 14833 -12011 14867
rect -11973 14833 -11939 14867
rect -11901 14833 -11867 14867
rect -11829 14833 -11795 14867
rect -11757 14833 -11723 14867
rect -11685 14833 -11651 14867
rect -11613 14833 -11579 14867
rect -11541 14833 -11507 14867
rect -11469 14833 -11435 14867
rect -11397 14833 -11363 14867
rect -11325 14833 -11291 14867
rect -11253 14833 -11219 14867
rect -11181 14833 -11147 14867
rect -11109 14833 -11075 14867
rect -11037 14833 -11003 14867
rect -10965 14833 -10931 14867
rect -10893 14833 -10859 14867
rect -10821 14833 -10787 14867
rect -10749 14833 -10715 14867
rect -10677 14833 -10643 14867
rect -10605 14833 -10571 14867
rect -10533 14833 -10499 14867
rect -10461 14833 -10427 14867
rect -10389 14833 -10355 14867
rect -10317 14833 -10283 14867
rect -10245 14833 -10211 14867
rect -10173 14833 -10139 14867
rect -10101 14833 -10067 14867
rect -10029 14833 -9995 14867
rect -9957 14833 -9923 14867
rect -9885 14833 -9851 14867
rect -9813 14833 -9779 14867
rect -9741 14833 -9707 14867
rect -9669 14833 -9635 14867
rect -9597 14833 -9563 14867
rect -9525 14833 -9491 14867
rect -9453 14833 -9419 14867
rect -9381 14833 -9347 14867
rect -9309 14833 -9275 14867
rect -9237 14833 -9203 14867
rect -9165 14833 -9131 14867
rect -9093 14833 -9059 14867
rect -9021 14833 -8987 14867
rect -8949 14833 -8915 14867
rect -8877 14833 -8843 14867
rect -8805 14833 -8771 14867
rect -8733 14833 -8699 14867
rect -8661 14833 -8627 14867
rect -8589 14833 -8555 14867
rect -8517 14833 -8483 14867
rect -8445 14833 -8411 14867
rect -8373 14833 -8339 14867
rect -8301 14833 -8267 14867
rect -8229 14833 -8195 14867
rect -8157 14833 -8123 14867
rect -8085 14833 -8051 14867
rect -8013 14833 -7979 14867
rect -7941 14833 -7907 14867
rect -7869 14833 -7835 14867
rect -7797 14833 -7763 14867
rect -7725 14833 -7691 14867
rect -7653 14833 -7619 14867
rect -7581 14833 -7547 14867
rect -7509 14833 -7475 14867
rect -7437 14833 -7403 14867
rect -7365 14833 -7331 14867
rect -7293 14833 -7259 14867
rect -7221 14833 -7187 14867
rect -7149 14833 -7115 14867
rect -7077 14833 -7043 14867
rect -7005 14833 -6971 14867
rect -6933 14833 -6899 14867
rect -6861 14833 -6827 14867
rect -6789 14833 -6755 14867
rect -6717 14833 -6683 14867
rect -6645 14833 -6611 14867
rect -6573 14833 -6539 14867
rect -6501 14833 -6467 14867
rect -6429 14833 -6395 14867
rect -6357 14833 -6323 14867
rect -6285 14833 -6251 14867
rect -6213 14833 -6179 14867
rect -6141 14833 -6107 14867
rect -6069 14833 -6035 14867
rect -5997 14833 -5963 14867
rect -5925 14833 -5891 14867
rect -5853 14833 -5819 14867
rect -5781 14833 -5747 14867
rect -5709 14833 -5675 14867
rect -5637 14833 -5603 14867
rect -5565 14833 -5531 14867
rect -5493 14833 -5459 14867
rect -5421 14833 -5387 14867
rect -5349 14833 -5315 14867
rect -5277 14833 -5243 14867
rect -5205 14833 -5171 14867
rect -5133 14833 -5099 14867
rect -5061 14833 -5027 14867
rect -4989 14833 -4955 14867
rect -4917 14833 -4883 14867
rect -4845 14833 -4811 14867
rect -4773 14833 -4739 14867
rect -4701 14833 -4667 14867
rect -4629 14833 -4595 14867
rect -4557 14833 -4523 14867
rect -4485 14833 -4451 14867
rect -4413 14833 -4379 14867
rect -4341 14833 -4307 14867
rect -4269 14833 -4235 14867
rect -4197 14833 -4163 14867
rect -4125 14833 -4091 14867
rect -4053 14833 -4019 14867
rect -3981 14833 -3947 14867
rect -3909 14833 -3875 14867
rect -3837 14833 -3803 14867
rect -3765 14833 -3731 14867
rect -3693 14833 -3659 14867
rect -3621 14833 -3587 14867
rect -3549 14833 -3515 14867
rect -3477 14833 -3443 14867
rect -3405 14833 -3371 14867
rect -3333 14833 -3299 14867
rect -3261 14833 -3227 14867
rect -3189 14833 -3155 14867
rect -3117 14833 -3083 14867
rect -3045 14833 -3011 14867
rect -2973 14833 -2939 14867
rect -2901 14833 -2867 14867
rect -2829 14833 -2795 14867
rect -2757 14833 -2723 14867
rect -2685 14833 -2651 14867
rect -2613 14833 -2579 14867
rect -2541 14833 -2507 14867
rect -2469 14833 -2435 14867
rect -2397 14833 -2363 14867
rect -2325 14833 -2291 14867
rect -2253 14833 -2219 14867
rect -2181 14833 -2147 14867
rect -2109 14833 -2075 14867
rect -2037 14833 -2003 14867
rect -1965 14833 -1931 14867
rect -1893 14833 -1859 14867
rect -1821 14833 -1787 14867
rect -1749 14833 -1715 14867
rect -1677 14833 -1643 14867
rect -1605 14833 -1571 14867
rect -1533 14833 -1499 14867
rect -1461 14833 -1427 14867
rect -1389 14833 -1355 14867
rect -1317 14833 -1283 14867
rect -1245 14833 -1211 14867
rect -1173 14833 -1139 14867
rect -1101 14833 -1067 14867
rect -1029 14833 -995 14867
rect -957 14833 -923 14867
rect -885 14833 -851 14867
rect -813 14833 -779 14867
rect -741 14833 -707 14867
rect -669 14833 -635 14867
rect -597 14833 -563 14867
rect -525 14833 -491 14867
rect -453 14833 -419 14867
rect -381 14833 -347 14867
rect -309 14833 -275 14867
rect -237 14833 -203 14867
rect -165 14833 -131 14867
rect -93 14833 -59 14867
rect -21 14833 13 14867
rect 51 14833 85 14867
rect 123 14833 157 14867
rect 195 14833 229 14867
rect 267 14833 301 14867
rect 339 14833 373 14867
rect 411 14833 445 14867
rect 483 14833 517 14867
rect 555 14833 589 14867
rect 627 14833 661 14867
rect 699 14833 733 14867
rect 771 14833 805 14867
rect 843 14833 877 14867
rect 915 14833 949 14867
rect 987 14833 1021 14867
rect 1059 14833 1093 14867
rect 1131 14833 1165 14867
rect 1203 14833 1237 14867
rect 1275 14833 1309 14867
rect 1347 14833 1381 14867
rect 1419 14833 1453 14867
rect 1491 14833 1525 14867
rect 1563 14833 1597 14867
rect 1635 14833 1669 14867
rect 1707 14833 1741 14867
rect 1779 14833 1813 14867
rect 1851 14833 1885 14867
rect 1923 14833 1957 14867
rect 1995 14833 2029 14867
rect 2067 14833 2101 14867
rect 2139 14833 2173 14867
rect 2211 14833 2245 14867
rect 2283 14833 2317 14867
rect 2355 14833 2389 14867
rect 2427 14833 2461 14867
rect 2499 14833 2533 14867
rect 2571 14833 2605 14867
rect 2643 14833 2677 14867
rect 2715 14833 2749 14867
rect 2787 14833 2821 14867
rect 2859 14833 2893 14867
rect 2931 14833 2965 14867
rect 3003 14833 3037 14867
rect 3075 14833 3109 14867
rect 3147 14833 3181 14867
rect 3219 14833 3253 14867
rect 3291 14833 3325 14867
rect 3363 14833 3397 14867
rect 3435 14833 3469 14867
rect 3507 14833 3541 14867
rect 3579 14833 3613 14867
rect 3651 14833 3685 14867
rect 3723 14833 3757 14867
rect 3795 14833 3829 14867
rect 3867 14833 3901 14867
rect 3939 14833 3973 14867
rect 4011 14833 4045 14867
rect 4083 14833 4117 14867
rect 4155 14833 4189 14867
rect 4227 14833 4261 14867
rect 4299 14833 4333 14867
rect 4371 14833 4405 14867
rect 4443 14833 4477 14867
rect 4515 14833 4549 14867
rect 4587 14833 4621 14867
rect 4659 14833 4693 14867
rect 4731 14833 4765 14867
rect 4803 14833 4837 14867
rect 4875 14833 4909 14867
rect 4947 14833 4981 14867
rect 5019 14833 5053 14867
rect 5091 14833 5125 14867
rect 5163 14833 5197 14867
rect 5235 14833 5269 14867
rect 5307 14833 5341 14867
rect 5379 14833 5413 14867
rect 5451 14833 5485 14867
rect 5523 14833 5557 14867
rect 5595 14833 5629 14867
rect 5667 14833 5701 14867
rect 5739 14833 5773 14867
rect 5811 14833 5845 14867
rect 5883 14833 5917 14867
rect 5955 14833 5989 14867
rect 6027 14833 6061 14867
rect 6099 14833 6133 14867
rect 6171 14833 6205 14867
rect 6243 14833 6277 14867
rect 6315 14833 6349 14867
rect 6387 14833 6421 14867
rect 6459 14833 6493 14867
rect 6531 14833 6565 14867
rect 6603 14833 6637 14867
rect 6675 14833 6709 14867
rect 6747 14833 6781 14867
rect 6819 14833 6853 14867
rect 6891 14833 6925 14867
rect 6963 14833 6997 14867
rect 7035 14833 7069 14867
rect 7107 14833 7141 14867
rect 7179 14833 7213 14867
rect 7251 14833 7285 14867
rect 7323 14833 7357 14867
rect 7395 14833 7429 14867
rect 7467 14833 7501 14867
rect 7539 14833 7573 14867
rect 7611 14833 7645 14867
rect 7683 14833 7717 14867
rect 7755 14833 7789 14867
rect 7827 14833 7861 14867
rect 7899 14833 7933 14867
rect 7971 14833 8005 14867
rect 8043 14833 8077 14867
rect 8115 14833 8149 14867
rect 8187 14833 8221 14867
rect 8259 14833 8293 14867
rect 8331 14833 8365 14867
rect 8403 14833 8437 14867
rect 8475 14833 8509 14867
rect 8547 14833 8581 14867
rect 8619 14833 8653 14867
rect 8691 14833 8725 14867
rect 8763 14833 8797 14867
rect 8835 14833 8869 14867
rect 8907 14833 8941 14867
rect 8979 14833 9013 14867
rect 9051 14833 9085 14867
rect 9123 14833 9157 14867
rect 9195 14833 9229 14867
rect 9267 14833 9301 14867
rect 9339 14833 9373 14867
rect 9411 14833 9445 14867
rect 9483 14833 9517 14867
rect 9555 14833 9589 14867
rect 9627 14833 9661 14867
rect 9699 14833 9733 14867
rect 9771 14833 9805 14867
rect 9843 14833 9877 14867
rect 9915 14833 9949 14867
rect 9987 14833 10021 14867
rect 10059 14833 10093 14867
rect 10131 14833 10165 14867
rect 10203 14833 10237 14867
rect 10275 14833 10309 14867
rect 10347 14833 10381 14867
rect 10419 14833 10453 14867
rect 10491 14833 10525 14867
rect 10563 14833 10597 14867
rect 10635 14833 10669 14867
rect 10707 14833 10741 14867
rect 10779 14833 10813 14867
rect 10851 14833 10885 14867
rect 10923 14833 10957 14867
rect 10995 14833 11029 14867
rect 11067 14833 11101 14867
rect 11139 14833 11173 14867
rect 11211 14833 11245 14867
rect 11283 14833 11317 14867
rect 11355 14833 11389 14867
rect 11427 14833 11461 14867
rect 11499 14833 11533 14867
rect 11571 14833 11605 14867
rect 11643 14833 11677 14867
rect 11715 14833 11749 14867
rect 11787 14833 11821 14867
rect 11859 14833 11893 14867
rect 11931 14833 11965 14867
rect 12003 14833 12037 14867
rect 12075 14833 12109 14867
rect 12147 14833 12181 14867
rect 12219 14833 12253 14867
rect 12291 14833 12325 14867
rect 12363 14833 12397 14867
rect 12435 14833 12469 14867
rect 12507 14833 12541 14867
rect 12579 14833 12613 14867
rect 12651 14833 12685 14867
rect 12723 14833 12757 14867
rect 12795 14833 12829 14867
rect 12867 14833 12901 14867
rect 12939 14833 12973 14867
rect 13011 14833 13045 14867
rect 13083 14833 13117 14867
rect 13155 14833 13189 14867
rect 13227 14833 13261 14867
rect 13299 14833 13333 14867
rect 13371 14833 13405 14867
rect 13443 14833 13477 14867
rect 13515 14833 13549 14867
rect 13587 14833 13621 14867
rect 13659 14833 13693 14867
rect 13731 14833 13765 14867
rect 13803 14833 13837 14867
rect 13875 14833 13909 14867
rect 13947 14833 13981 14867
rect 14019 14833 14053 14867
rect 14091 14833 14125 14867
rect 14163 14833 14197 14867
rect 14235 14833 14269 14867
rect 14307 14833 14341 14867
rect 14379 14833 14413 14867
rect 14451 14833 14485 14867
rect 14523 14833 14557 14867
rect 14595 14833 14629 14867
rect 14667 14833 14701 14867
rect 14739 14833 14773 14867
rect 14811 14833 14845 14867
rect 14883 14833 14917 14867
rect 14955 14833 14989 14867
rect 15027 14833 15061 14867
rect 15099 14833 15133 14867
rect 15171 14833 15205 14867
rect 15243 14833 15277 14867
rect 15315 14833 15349 14867
rect 15387 14833 15421 14867
rect 15459 14833 15493 14867
rect 15531 14833 15565 14867
rect 15603 14833 15637 14867
rect 15675 14833 15709 14867
rect 15747 14833 15781 14867
rect 15819 14833 15853 14867
rect 15891 14833 15925 14867
rect 15963 14833 15997 14867
rect 16035 14833 16069 14867
rect 16107 14833 16141 14867
rect 16179 14833 16213 14867
rect 16251 14833 16285 14867
rect 16323 14833 16357 14867
rect 16395 14833 16429 14867
rect 16467 14833 16501 14867
rect 16539 14833 16573 14867
rect 16611 14833 16645 14867
rect 16683 14833 16717 14867
rect 16755 14833 16789 14867
rect 16827 14833 16861 14867
rect 16899 14833 16933 14867
rect 16971 14833 17005 14867
rect 17043 14833 17077 14867
rect 17115 14833 17149 14867
rect 17187 14833 17221 14867
rect 17259 14833 17293 14867
rect 17331 14833 17365 14867
rect 17403 14833 17437 14867
rect 17475 14833 17509 14867
rect 17547 14833 17581 14867
rect 17619 14833 17653 14867
rect 17691 14833 17725 14867
rect 17763 14833 17797 14867
rect 17835 14833 17869 14867
rect 17907 14833 17941 14867
rect 17979 14833 18013 14867
rect 18051 14833 18085 14867
rect 18123 14833 18157 14867
rect 18195 14833 18229 14867
rect 18267 14833 18301 14867
rect 18339 14833 18373 14867
rect 18411 14833 18445 14867
rect 18483 14833 18517 14867
rect 18555 14833 18589 14867
rect 18627 14833 18661 14867
rect 18699 14833 18733 14867
rect 18771 14833 18805 14867
rect 18843 14833 18877 14867
rect 18915 14833 18949 14867
rect 18987 14833 19021 14867
rect 19059 14833 19093 14867
rect 19131 14833 19165 14867
rect 19203 14833 19237 14867
rect 19275 14833 19309 14867
rect 19347 14833 19381 14867
rect 19419 14833 19453 14867
rect 19491 14833 19525 14867
rect 19563 14833 19597 14867
rect 19635 14833 19669 14867
rect 19707 14833 19741 14867
rect 19779 14833 19813 14867
rect 19851 14833 19885 14867
rect 19923 14833 19957 14867
rect 19995 14833 20029 14867
rect 20067 14833 20101 14867
rect 20139 14833 20173 14867
rect 20211 14833 20245 14867
rect 20283 14833 20317 14867
rect 20355 14833 20389 14867
rect 20427 14833 20461 14867
rect 20499 14833 20533 14867
rect 20571 14833 20605 14867
rect 20643 14833 20677 14867
rect 20715 14833 20749 14867
rect 20787 14833 20821 14867
rect 20859 14833 20893 14867
rect 20931 14833 20965 14867
rect 21003 14833 21037 14867
rect 21075 14833 21109 14867
rect 21147 14833 21181 14867
rect 21219 14833 21253 14867
rect 21291 14833 21325 14867
rect 21363 14833 21397 14867
rect 21435 14833 21469 14867
rect 21507 14833 21541 14867
rect 21579 14833 21613 14867
rect 21651 14833 21685 14867
rect 21723 14833 21757 14867
rect 21795 14833 21829 14867
rect 21867 14833 21901 14867
rect 21939 14833 21973 14867
rect 22011 14833 22045 14867
rect 22083 14833 22117 14867
rect 22155 14833 22189 14867
rect 22227 14833 22261 14867
rect 22299 14833 22333 14867
rect 22371 14833 22405 14867
rect 22443 14833 22477 14867
rect 22515 14833 22549 14867
rect 22587 14833 22621 14867
rect 22659 14833 22693 14867
rect 22731 14833 22765 14867
rect 22803 14833 22837 14867
rect 22875 14833 22909 14867
rect 22947 14833 22981 14867
rect 23019 14833 23053 14867
rect 23091 14833 23125 14867
rect 23163 14833 23197 14867
rect 23235 14833 23269 14867
rect 23307 14833 23341 14867
rect 23379 14833 23413 14867
rect 23451 14833 23485 14867
rect 23523 14833 23557 14867
rect 23595 14833 23629 14867
rect 23667 14833 23701 14867
rect 23739 14833 23773 14867
rect 23811 14833 23845 14867
rect 23883 14833 23917 14867
rect 23955 14833 23989 14867
rect 24027 14833 24061 14867
rect 24099 14833 24133 14867
rect 24171 14833 24205 14867
rect 24243 14833 24277 14867
rect 24315 14833 24349 14867
rect 24387 14833 24421 14867
rect 24459 14833 24493 14867
rect 24531 14833 24565 14867
rect 24603 14833 24637 14867
rect 24675 14833 24709 14867
rect 24747 14833 24781 14867
rect 24819 14833 24853 14867
rect 24891 14833 24925 14867
rect 24963 14833 24997 14867
rect 25035 14833 25069 14867
rect 25107 14833 25141 14867
rect 25179 14833 25213 14867
rect 25251 14833 25285 14867
rect 25323 14833 25357 14867
rect 25395 14833 25429 14867
rect 25467 14833 25501 14867
rect 25539 14833 25573 14867
rect 25611 14833 25645 14867
rect 25683 14833 25717 14867
rect 25755 14833 25789 14867
rect 25827 14833 25861 14867
rect 25899 14833 25933 14867
rect 25971 14833 26005 14867
rect 26043 14833 26077 14867
rect 26115 14833 26149 14867
rect 26187 14833 26221 14867
rect 26259 14833 26293 14867
rect 26331 14833 26365 14867
rect 26403 14833 26437 14867
rect 26475 14833 26509 14867
rect 26547 14833 26581 14867
rect 26619 14833 26653 14867
rect 26691 14833 26725 14867
rect 26763 14833 26797 14867
rect 26835 14833 26869 14867
rect 26907 14833 26941 14867
rect 26979 14833 27013 14867
rect 27051 14833 27085 14867
rect 27123 14833 27157 14867
rect 27195 14833 27229 14867
rect 27267 14833 27301 14867
rect 27339 14833 27373 14867
rect 27411 14833 27445 14867
rect 27483 14833 27517 14867
rect 27555 14833 27589 14867
rect 27627 14833 27661 14867
rect 27699 14833 27733 14867
rect 27771 14833 27805 14867
rect 27843 14833 27877 14867
rect 27915 14833 27949 14867
rect 27987 14833 28021 14867
rect 28059 14833 28093 14867
rect 28131 14833 28165 14867
rect 28203 14833 28237 14867
rect 28275 14833 28309 14867
rect 28347 14833 28381 14867
rect 28419 14833 28453 14867
rect 28491 14833 28525 14867
rect 28563 14833 28597 14867
rect 28635 14833 28669 14867
rect 28707 14833 28741 14867
rect 28779 14833 28813 14867
rect 28851 14833 28885 14867
rect 28923 14833 28957 14867
rect 28995 14833 29029 14867
rect 29067 14833 29101 14867
rect 29139 14833 29173 14867
rect 29211 14833 29245 14867
rect 29283 14833 29317 14867
rect 29355 14833 29389 14867
rect 29427 14833 29461 14867
rect 29499 14833 29533 14867
rect 29571 14833 29605 14867
rect 29643 14833 29677 14867
rect 29715 14833 29749 14867
rect 29787 14833 29821 14867
rect 29859 14833 29893 14867
rect 29931 14833 29965 14867
rect 30003 14833 30037 14867
rect 30075 14833 30109 14867
rect 30147 14833 30181 14867
rect 30219 14833 30253 14867
rect 30291 14833 30325 14867
rect 30363 14833 30397 14867
rect 30435 14833 30469 14867
rect 30507 14833 30541 14867
rect 30579 14833 30613 14867
rect 30651 14833 30685 14867
rect 30723 14833 30757 14867
rect 30795 14833 30829 14867
rect 30867 14833 30901 14867
rect 30939 14833 30973 14867
rect 31011 14833 31045 14867
rect 31083 14833 31117 14867
rect 31155 14833 31189 14867
rect 31227 14833 31261 14867
rect 31299 14833 31333 14867
rect 31371 14833 31405 14867
rect 31443 14833 31477 14867
rect 31515 14833 31549 14867
rect 31587 14833 31621 14867
rect 31659 14833 31693 14867
rect 31731 14833 31765 14867
rect 31803 14833 31837 14867
rect 31875 14833 31909 14867
rect 31947 14833 31981 14867
rect 32019 14833 32053 14867
rect 32091 14833 32125 14867
rect 32163 14833 32197 14867
rect 32235 14833 32269 14867
rect 32307 14833 32341 14867
rect 32379 14833 32413 14867
rect 32451 14833 32485 14867
rect 32523 14833 32557 14867
rect 32595 14833 32629 14867
rect 32667 14833 32701 14867
rect 32739 14833 32773 14867
rect 32811 14833 32845 14867
rect 32883 14833 32917 14867
rect 32955 14833 32989 14867
rect 33027 14833 33061 14867
rect 33099 14833 33133 14867
rect 33171 14833 33205 14867
rect 33243 14833 33277 14867
rect 33315 14833 33349 14867
rect 33387 14833 33421 14867
rect 33459 14833 33493 14867
rect 33531 14833 33565 14867
rect 33603 14833 33637 14867
rect 33675 14833 33709 14867
rect 33747 14833 33781 14867
rect 33819 14833 33853 14867
rect 33891 14833 33925 14867
rect 33963 14833 33997 14867
rect 34035 14833 34069 14867
rect 34107 14833 34141 14867
rect 34179 14833 34213 14867
rect 34251 14833 34285 14867
rect 34323 14833 34357 14867
rect 34395 14833 34429 14867
rect 34467 14833 34501 14867
rect 34539 14833 34573 14867
rect 34611 14833 34645 14867
rect 34683 14833 34717 14867
rect 34755 14833 34789 14867
rect 34827 14833 34861 14867
rect 34899 14833 34933 14867
rect 34971 14833 35005 14867
rect 35043 14833 35077 14867
rect 35115 14833 35149 14867
rect 35187 14833 35221 14867
rect -17467 14763 -17433 14797
rect -17467 14691 -17433 14725
rect -17467 14619 -17433 14653
rect -17467 14547 -17433 14581
rect -17467 14475 -17433 14509
rect -17467 14403 -17433 14437
rect -17467 14331 -17433 14365
rect -17467 14259 -17433 14293
rect -17467 14187 -17433 14221
rect -17467 14115 -17433 14149
rect -17467 14043 -17433 14077
rect -17467 13971 -17433 14005
rect -17467 13899 -17433 13933
rect 35333 14763 35367 14797
rect 35333 14691 35367 14725
rect 35333 14619 35367 14653
rect 35333 14547 35367 14581
rect 35333 14475 35367 14509
rect 35333 14403 35367 14437
rect 35333 14331 35367 14365
rect 35333 14259 35367 14293
rect 35333 14187 35367 14221
rect 35333 14115 35367 14149
rect 35333 14043 35367 14077
rect 35333 13971 35367 14005
rect 35333 13899 35367 13933
rect -17467 13827 -17433 13861
rect -17467 13755 -17433 13789
rect -17467 13683 -17433 13717
rect -17467 13611 -17433 13645
rect -17467 13539 -17433 13573
rect -17467 13467 -17433 13501
rect -17467 13395 -17433 13429
rect -17467 13323 -17433 13357
rect -17467 13251 -17433 13285
rect -17467 13179 -17433 13213
rect -17467 13107 -17433 13141
rect -17467 13035 -17433 13069
rect -17467 12963 -17433 12997
rect -17467 12891 -17433 12925
rect -17467 12819 -17433 12853
rect -17467 12747 -17433 12781
rect -17467 12675 -17433 12709
rect -17467 12603 -17433 12637
rect -17467 12531 -17433 12565
rect -17467 12459 -17433 12493
rect -17467 12387 -17433 12421
rect -17467 12315 -17433 12349
rect -17467 12243 -17433 12277
rect -17467 12171 -17433 12205
rect -17467 12099 -17433 12133
rect 35333 13827 35367 13861
rect 35333 13755 35367 13789
rect 35333 13683 35367 13717
rect 35333 13611 35367 13645
rect 35333 13539 35367 13573
rect 35333 13467 35367 13501
rect 35333 13395 35367 13429
rect 35333 13323 35367 13357
rect 35333 13251 35367 13285
rect 35333 13179 35367 13213
rect 35333 13107 35367 13141
rect 35333 13035 35367 13069
rect 35333 12963 35367 12997
rect 35333 12891 35367 12925
rect 35333 12819 35367 12853
rect 35333 12747 35367 12781
rect 35333 12675 35367 12709
rect 35333 12603 35367 12637
rect 35333 12531 35367 12565
rect 35333 12459 35367 12493
rect 35333 12387 35367 12421
rect 35333 12315 35367 12349
rect 35333 12243 35367 12277
rect 35333 12171 35367 12205
rect 35333 12099 35367 12133
rect -17467 12027 -17433 12061
rect -17467 11955 -17433 11989
rect -17467 11883 -17433 11917
rect -17467 11811 -17433 11845
rect -17467 11739 -17433 11773
rect -17467 11667 -17433 11701
rect -17467 11595 -17433 11629
rect -17467 11523 -17433 11557
rect -17467 11451 -17433 11485
rect -17467 11379 -17433 11413
rect -17467 11307 -17433 11341
rect -17467 11235 -17433 11269
rect -17467 11163 -17433 11197
rect -17467 11091 -17433 11125
rect -17467 11019 -17433 11053
rect -17467 10947 -17433 10981
rect -17467 10875 -17433 10909
rect -17467 10803 -17433 10837
rect -17467 10731 -17433 10765
rect -17467 10659 -17433 10693
rect -17467 10587 -17433 10621
rect -17467 10515 -17433 10549
rect -17467 10443 -17433 10477
rect 35333 12027 35367 12061
rect 35333 11955 35367 11989
rect 35333 11883 35367 11917
rect 35333 11811 35367 11845
rect 35333 11739 35367 11773
rect 35333 11667 35367 11701
rect 35333 11595 35367 11629
rect 35333 11523 35367 11557
rect 35333 11451 35367 11485
rect 35333 11379 35367 11413
rect 35333 11307 35367 11341
rect 35333 11235 35367 11269
rect 35333 11163 35367 11197
rect 35333 11091 35367 11125
rect 35333 11019 35367 11053
rect 35333 10947 35367 10981
rect 35333 10875 35367 10909
rect 35333 10803 35367 10837
rect 35333 10731 35367 10765
rect 35333 10659 35367 10693
rect 35333 10587 35367 10621
rect 35333 10515 35367 10549
rect 35333 10443 35367 10477
rect -17467 10371 -17433 10405
rect 35333 10371 35367 10405
rect -17467 10299 -17433 10333
rect -17467 10227 -17433 10261
rect -17467 10155 -17433 10189
rect -17467 10083 -17433 10117
rect -17467 10011 -17433 10045
rect -17467 9939 -17433 9973
rect -17467 9867 -17433 9901
rect -17467 9795 -17433 9829
rect -17467 9723 -17433 9757
rect -17467 9651 -17433 9685
rect -17467 9579 -17433 9613
rect -17467 9507 -17433 9541
rect -17467 9435 -17433 9469
rect -17467 9363 -17433 9397
rect -17467 9291 -17433 9325
rect -17467 9219 -17433 9253
rect -17467 9147 -17433 9181
rect -17467 9075 -17433 9109
rect -17467 9003 -17433 9037
rect -17467 8931 -17433 8965
rect -17467 8859 -17433 8893
rect -17467 8787 -17433 8821
rect -17467 8715 -17433 8749
rect -17467 8643 -17433 8677
rect -17467 8571 -17433 8605
rect 35333 10299 35367 10333
rect 35333 10227 35367 10261
rect 35333 10155 35367 10189
rect 35333 10083 35367 10117
rect 35333 10011 35367 10045
rect 35333 9939 35367 9973
rect 35333 9867 35367 9901
rect 35333 9795 35367 9829
rect 35333 9723 35367 9757
rect 35333 9651 35367 9685
rect 35333 9579 35367 9613
rect 35333 9507 35367 9541
rect 35333 9435 35367 9469
rect 35333 9363 35367 9397
rect 35333 9291 35367 9325
rect 35333 9219 35367 9253
rect 35333 9147 35367 9181
rect 35333 9075 35367 9109
rect 35333 9003 35367 9037
rect 35333 8931 35367 8965
rect 35333 8859 35367 8893
rect 35333 8787 35367 8821
rect 35333 8715 35367 8749
rect 35333 8643 35367 8677
rect 35333 8571 35367 8605
rect -17467 8499 -17433 8533
rect -17467 8427 -17433 8461
rect -17467 8355 -17433 8389
rect -17467 8283 -17433 8317
rect -17467 8211 -17433 8245
rect -17467 8139 -17433 8173
rect -17467 8067 -17433 8101
rect -17467 7995 -17433 8029
rect -17467 7923 -17433 7957
rect -17467 7851 -17433 7885
rect -17467 7779 -17433 7813
rect -17467 7707 -17433 7741
rect -17467 7635 -17433 7669
rect -17467 7563 -17433 7597
rect -17467 7491 -17433 7525
rect -17467 7419 -17433 7453
rect -17467 7347 -17433 7381
rect -17467 7275 -17433 7309
rect -17467 7203 -17433 7237
rect -17467 7131 -17433 7165
rect -17467 7059 -17433 7093
rect -17467 6987 -17433 7021
rect -17467 6915 -17433 6949
rect -17467 6843 -17433 6877
rect -17467 6771 -17433 6805
rect -17467 6699 -17433 6733
rect -17467 6627 -17433 6661
rect -17467 6555 -17433 6589
rect 35333 8499 35367 8533
rect 35333 8427 35367 8461
rect 35333 8355 35367 8389
rect 35333 8283 35367 8317
rect 35333 8211 35367 8245
rect 35333 8139 35367 8173
rect 35333 8067 35367 8101
rect 35333 7995 35367 8029
rect 35333 7923 35367 7957
rect 35333 7851 35367 7885
rect 35333 7779 35367 7813
rect 35333 7707 35367 7741
rect 35333 7635 35367 7669
rect 35333 7563 35367 7597
rect 35333 7491 35367 7525
rect 35333 7419 35367 7453
rect 35333 7347 35367 7381
rect 35333 7275 35367 7309
rect 35333 7203 35367 7237
rect 35333 7131 35367 7165
rect 35333 7059 35367 7093
rect 35333 6987 35367 7021
rect 35333 6915 35367 6949
rect 35333 6843 35367 6877
rect 35333 6771 35367 6805
rect 35333 6699 35367 6733
rect 35333 6627 35367 6661
rect 35333 6555 35367 6589
rect -17467 6483 -17433 6517
rect 35333 6483 35367 6517
rect -17467 6411 -17433 6445
rect -17467 6339 -17433 6373
rect -17467 6267 -17433 6301
rect -17467 6195 -17433 6229
rect -17467 6123 -17433 6157
rect -17467 6051 -17433 6085
rect -17467 5979 -17433 6013
rect -17467 5907 -17433 5941
rect -17467 5835 -17433 5869
rect -17467 5763 -17433 5797
rect -17467 5691 -17433 5725
rect -17467 5619 -17433 5653
rect -17467 5547 -17433 5581
rect -17467 5475 -17433 5509
rect -17467 5403 -17433 5437
rect -17467 5331 -17433 5365
rect -17467 5259 -17433 5293
rect -17467 5187 -17433 5221
rect -17467 5115 -17433 5149
rect -17467 5043 -17433 5077
rect -17467 4971 -17433 5005
rect -17467 4899 -17433 4933
rect -17467 4827 -17433 4861
rect -17467 4755 -17433 4789
rect -17467 4683 -17433 4717
rect 35333 6411 35367 6445
rect 35333 6339 35367 6373
rect 35333 6267 35367 6301
rect 35333 6195 35367 6229
rect 35333 6123 35367 6157
rect 35333 6051 35367 6085
rect 35333 5979 35367 6013
rect 35333 5907 35367 5941
rect 35333 5835 35367 5869
rect 35333 5763 35367 5797
rect 35333 5691 35367 5725
rect 35333 5619 35367 5653
rect 35333 5547 35367 5581
rect 35333 5475 35367 5509
rect 35333 5403 35367 5437
rect 35333 5331 35367 5365
rect 35333 5259 35367 5293
rect 35333 5187 35367 5221
rect 35333 5115 35367 5149
rect 35333 5043 35367 5077
rect 35333 4971 35367 5005
rect 35333 4899 35367 4933
rect 35333 4827 35367 4861
rect 35333 4755 35367 4789
rect -17467 4611 -17433 4645
rect 35333 4683 35367 4717
rect -17467 4539 -17433 4573
rect -17467 4467 -17433 4501
rect -17467 4395 -17433 4429
rect -17467 4323 -17433 4357
rect -17467 4251 -17433 4285
rect -17467 4179 -17433 4213
rect -17467 4107 -17433 4141
rect -17467 4035 -17433 4069
rect -17467 3963 -17433 3997
rect -17467 3891 -17433 3925
rect -17467 3819 -17433 3853
rect -17467 3747 -17433 3781
rect -17467 3675 -17433 3709
rect -17467 3603 -17433 3637
rect -17467 3531 -17433 3565
rect -17467 3459 -17433 3493
rect -17467 3387 -17433 3421
rect -17467 3315 -17433 3349
rect -17467 3243 -17433 3277
rect -17467 3171 -17433 3205
rect -17467 3099 -17433 3133
rect -17467 3027 -17433 3061
rect 35333 4611 35367 4645
rect 35333 4539 35367 4573
rect 35333 4467 35367 4501
rect 35333 4395 35367 4429
rect 35333 4323 35367 4357
rect 35333 4251 35367 4285
rect 35333 4179 35367 4213
rect 35333 4107 35367 4141
rect 35333 4035 35367 4069
rect 35333 3963 35367 3997
rect 35333 3891 35367 3925
rect 35333 3819 35367 3853
rect 35333 3747 35367 3781
rect 35333 3675 35367 3709
rect 35333 3603 35367 3637
rect 35333 3531 35367 3565
rect 35333 3459 35367 3493
rect 35333 3387 35367 3421
rect 35333 3315 35367 3349
rect 35333 3243 35367 3277
rect 35333 3171 35367 3205
rect 35333 3099 35367 3133
rect 35333 3027 35367 3061
rect -17467 2955 -17433 2989
rect -17467 2883 -17433 2917
rect -17467 2811 -17433 2845
rect -17467 2739 -17433 2773
rect -17467 2667 -17433 2701
rect -17467 2595 -17433 2629
rect -17467 2523 -17433 2557
rect -17467 2451 -17433 2485
rect -17467 2379 -17433 2413
rect -17467 2307 -17433 2341
rect -17467 2235 -17433 2269
rect -17467 2163 -17433 2197
rect -17467 2091 -17433 2125
rect -17467 2019 -17433 2053
rect -17467 1947 -17433 1981
rect -17467 1875 -17433 1909
rect -17467 1803 -17433 1837
rect -17467 1731 -17433 1765
rect -17467 1659 -17433 1693
rect -17467 1587 -17433 1621
rect -17467 1515 -17433 1549
rect -17467 1443 -17433 1477
rect -17467 1371 -17433 1405
rect -17467 1299 -17433 1333
rect -17467 1227 -17433 1261
rect 35333 2955 35367 2989
rect 35333 2883 35367 2917
rect 35333 2811 35367 2845
rect 35333 2739 35367 2773
rect 35333 2667 35367 2701
rect 35333 2595 35367 2629
rect 35333 2523 35367 2557
rect 35333 2451 35367 2485
rect 35333 2379 35367 2413
rect 35333 2307 35367 2341
rect 35333 2235 35367 2269
rect 35333 2163 35367 2197
rect 35333 2091 35367 2125
rect 35333 2019 35367 2053
rect 35333 1947 35367 1981
rect 35333 1875 35367 1909
rect 35333 1803 35367 1837
rect 35333 1731 35367 1765
rect 35333 1659 35367 1693
rect 35333 1587 35367 1621
rect 35333 1515 35367 1549
rect 35333 1443 35367 1477
rect 35333 1371 35367 1405
rect 35333 1299 35367 1333
rect 35333 1227 35367 1261
rect -17467 1155 -17433 1189
rect 35333 1155 35367 1189
rect -17467 1083 -17433 1117
rect -17467 1011 -17433 1045
rect -17467 939 -17433 973
rect -17467 867 -17433 901
rect -17467 795 -17433 829
rect -17467 723 -17433 757
rect -17467 651 -17433 685
rect -17467 579 -17433 613
rect -17467 507 -17433 541
rect -17467 435 -17433 469
rect -17467 363 -17433 397
rect -17467 291 -17433 325
rect -17467 219 -17433 253
rect -17467 147 -17433 181
rect -17467 75 -17433 109
rect -17467 3 -17433 37
rect -17467 -69 -17433 -35
rect -17467 -141 -17433 -107
rect -17467 -213 -17433 -179
rect -17467 -285 -17433 -251
rect -17467 -357 -17433 -323
rect -17467 -429 -17433 -395
rect -17467 -501 -17433 -467
rect -17467 -573 -17433 -539
rect -17467 -645 -17433 -611
rect -17467 -717 -17433 -683
rect -17467 -789 -17433 -755
rect -17467 -861 -17433 -827
rect 35333 1083 35367 1117
rect 35333 1011 35367 1045
rect 35333 939 35367 973
rect 35333 867 35367 901
rect 35333 795 35367 829
rect 35333 723 35367 757
rect 35333 651 35367 685
rect 35333 579 35367 613
rect 35333 507 35367 541
rect 35333 435 35367 469
rect 35333 363 35367 397
rect 35333 291 35367 325
rect 35333 219 35367 253
rect 35333 147 35367 181
rect 35333 75 35367 109
rect 35333 3 35367 37
rect 35333 -69 35367 -35
rect 35333 -141 35367 -107
rect 35333 -213 35367 -179
rect 35333 -285 35367 -251
rect 35333 -357 35367 -323
rect 35333 -429 35367 -395
rect 35333 -501 35367 -467
rect 35333 -573 35367 -539
rect 35333 -645 35367 -611
rect 35333 -717 35367 -683
rect 35333 -789 35367 -755
rect 35333 -861 35367 -827
rect -17467 -933 -17433 -899
rect 35333 -933 35367 -899
rect -17467 -1005 -17433 -971
rect -17467 -1077 -17433 -1043
rect -17467 -1149 -17433 -1115
rect -17467 -1221 -17433 -1187
rect -17467 -1293 -17433 -1259
rect -17467 -1365 -17433 -1331
rect -17467 -1437 -17433 -1403
rect -17467 -1509 -17433 -1475
rect -17467 -1581 -17433 -1547
rect -17467 -1653 -17433 -1619
rect -17467 -1725 -17433 -1691
rect -17467 -1797 -17433 -1763
rect -17467 -1869 -17433 -1835
rect -17467 -1941 -17433 -1907
rect -17467 -2013 -17433 -1979
rect -17467 -2085 -17433 -2051
rect -17467 -2157 -17433 -2123
rect -17467 -2229 -17433 -2195
rect -17467 -2301 -17433 -2267
rect -17467 -2373 -17433 -2339
rect -17467 -2445 -17433 -2411
rect -17467 -2517 -17433 -2483
rect -17467 -2589 -17433 -2555
rect -17467 -2661 -17433 -2627
rect -17467 -2733 -17433 -2699
rect 35333 -1005 35367 -971
rect 35333 -1077 35367 -1043
rect 35333 -1149 35367 -1115
rect 35333 -1221 35367 -1187
rect 35333 -1293 35367 -1259
rect 35333 -1365 35367 -1331
rect 35333 -1437 35367 -1403
rect 35333 -1509 35367 -1475
rect 35333 -1581 35367 -1547
rect 35333 -1653 35367 -1619
rect 35333 -1725 35367 -1691
rect 35333 -1797 35367 -1763
rect 35333 -1869 35367 -1835
rect 35333 -1941 35367 -1907
rect 35333 -2013 35367 -1979
rect 35333 -2085 35367 -2051
rect 35333 -2157 35367 -2123
rect 35333 -2229 35367 -2195
rect 35333 -2301 35367 -2267
rect 35333 -2373 35367 -2339
rect 35333 -2445 35367 -2411
rect 35333 -2517 35367 -2483
rect 35333 -2589 35367 -2555
rect 35333 -2661 35367 -2627
rect 35333 -2733 35367 -2699
rect -17467 -2805 -17433 -2771
rect -17467 -2877 -17433 -2843
rect -17467 -2949 -17433 -2915
rect -17467 -3021 -17433 -2987
rect -17467 -3093 -17433 -3059
rect -17467 -3165 -17433 -3131
rect -17467 -3237 -17433 -3203
rect -17467 -3309 -17433 -3275
rect -17467 -3381 -17433 -3347
rect -17467 -3453 -17433 -3419
rect -17467 -3525 -17433 -3491
rect -17467 -3597 -17433 -3563
rect -17467 -3669 -17433 -3635
rect -17467 -3741 -17433 -3707
rect -17467 -3813 -17433 -3779
rect -17467 -3885 -17433 -3851
rect -17467 -3957 -17433 -3923
rect -17467 -4029 -17433 -3995
rect -17467 -4101 -17433 -4067
rect -17467 -4173 -17433 -4139
rect -17467 -4245 -17433 -4211
rect -17467 -4317 -17433 -4283
rect -17467 -4389 -17433 -4355
rect 35333 -2805 35367 -2771
rect 35333 -2877 35367 -2843
rect 35333 -2949 35367 -2915
rect 35333 -3021 35367 -2987
rect 35333 -3093 35367 -3059
rect 35333 -3165 35367 -3131
rect 35333 -3237 35367 -3203
rect 35333 -3309 35367 -3275
rect 35333 -3381 35367 -3347
rect 35333 -3453 35367 -3419
rect 35333 -3525 35367 -3491
rect 35333 -3597 35367 -3563
rect 35333 -3669 35367 -3635
rect 35333 -3741 35367 -3707
rect 35333 -3813 35367 -3779
rect 35333 -3885 35367 -3851
rect 35333 -3957 35367 -3923
rect 35333 -4029 35367 -3995
rect 35333 -4101 35367 -4067
rect 35333 -4173 35367 -4139
rect 35333 -4245 35367 -4211
rect 35333 -4317 35367 -4283
rect 35333 -4389 35367 -4355
rect -17467 -4461 -17433 -4427
rect -17467 -4533 -17433 -4499
rect -17467 -4605 -17433 -4571
rect -17467 -4677 -17433 -4643
rect -17467 -4749 -17433 -4715
rect -17467 -4821 -17433 -4787
rect -17467 -4893 -17433 -4859
rect -17467 -4965 -17433 -4931
rect -17467 -5037 -17433 -5003
rect -17467 -5109 -17433 -5075
rect -17467 -5181 -17433 -5147
rect -17467 -5253 -17433 -5219
rect -17467 -5325 -17433 -5291
rect -17467 -5397 -17433 -5363
rect -17467 -5469 -17433 -5435
rect -17467 -5541 -17433 -5507
rect -17467 -5613 -17433 -5579
rect -17467 -5685 -17433 -5651
rect -17467 -5757 -17433 -5723
rect -17467 -5829 -17433 -5795
rect -17467 -5901 -17433 -5867
rect -17467 -5973 -17433 -5939
rect -17467 -6045 -17433 -6011
rect -17467 -6117 -17433 -6083
rect -17467 -6189 -17433 -6155
rect 35333 -4461 35367 -4427
rect 35333 -4533 35367 -4499
rect 35333 -4605 35367 -4571
rect 35333 -4677 35367 -4643
rect 35333 -4749 35367 -4715
rect 35333 -4821 35367 -4787
rect 35333 -4893 35367 -4859
rect 35333 -4965 35367 -4931
rect 35333 -5037 35367 -5003
rect 35333 -5109 35367 -5075
rect 35333 -5181 35367 -5147
rect 35333 -5253 35367 -5219
rect 35333 -5325 35367 -5291
rect 35333 -5397 35367 -5363
rect 35333 -5469 35367 -5435
rect 35333 -5541 35367 -5507
rect 35333 -5613 35367 -5579
rect 35333 -5685 35367 -5651
rect 35333 -5757 35367 -5723
rect 35333 -5829 35367 -5795
rect 35333 -5901 35367 -5867
rect 35333 -5973 35367 -5939
rect 35333 -6045 35367 -6011
rect 35333 -6117 35367 -6083
rect 35333 -6189 35367 -6155
rect -17467 -6261 -17433 -6227
rect -17467 -6333 -17433 -6299
rect -17467 -6405 -17433 -6371
rect -17467 -6477 -17433 -6443
rect -17467 -6549 -17433 -6515
rect -17467 -6621 -17433 -6587
rect -17467 -6693 -17433 -6659
rect -17467 -6765 -17433 -6731
rect -17467 -6837 -17433 -6803
rect -17467 -6909 -17433 -6875
rect -17467 -6981 -17433 -6947
rect -17467 -7053 -17433 -7019
rect -17467 -7125 -17433 -7091
rect -17467 -7197 -17433 -7163
rect 35333 -6261 35367 -6227
rect 35333 -6333 35367 -6299
rect 35333 -6405 35367 -6371
rect 35333 -6477 35367 -6443
rect 35333 -6549 35367 -6515
rect 35333 -6621 35367 -6587
rect 35333 -6693 35367 -6659
rect 35333 -6765 35367 -6731
rect 35333 -6837 35367 -6803
rect 35333 -6909 35367 -6875
rect 35333 -6981 35367 -6947
rect 35333 -7053 35367 -7019
rect 35333 -7125 35367 -7091
rect 35333 -7197 35367 -7163
rect -17321 -7267 -17287 -7233
rect -17249 -7267 -17215 -7233
rect -17177 -7267 -17143 -7233
rect -17105 -7267 -17071 -7233
rect -17033 -7267 -16999 -7233
rect -16961 -7267 -16927 -7233
rect -16889 -7267 -16855 -7233
rect -16817 -7267 -16783 -7233
rect -16745 -7267 -16711 -7233
rect -16673 -7267 -16639 -7233
rect -16601 -7267 -16567 -7233
rect -16529 -7267 -16495 -7233
rect -16457 -7267 -16423 -7233
rect -16385 -7267 -16351 -7233
rect -16313 -7267 -16279 -7233
rect -16241 -7267 -16207 -7233
rect -16169 -7267 -16135 -7233
rect -16097 -7267 -16063 -7233
rect -16025 -7267 -15991 -7233
rect -15953 -7267 -15919 -7233
rect -15881 -7267 -15847 -7233
rect -15809 -7267 -15775 -7233
rect -15737 -7267 -15703 -7233
rect -15665 -7267 -15631 -7233
rect -15593 -7267 -15559 -7233
rect -15521 -7267 -15487 -7233
rect -15449 -7267 -15415 -7233
rect -15377 -7267 -15343 -7233
rect -15305 -7267 -15271 -7233
rect -15233 -7267 -15199 -7233
rect -15161 -7267 -15127 -7233
rect -15089 -7267 -15055 -7233
rect -15017 -7267 -14983 -7233
rect -14945 -7267 -14911 -7233
rect -14873 -7267 -14839 -7233
rect -14801 -7267 -14767 -7233
rect -14729 -7267 -14695 -7233
rect -14657 -7267 -14623 -7233
rect -14585 -7267 -14551 -7233
rect -14513 -7267 -14479 -7233
rect -14441 -7267 -14407 -7233
rect -14369 -7267 -14335 -7233
rect -14297 -7267 -14263 -7233
rect -14225 -7267 -14191 -7233
rect -14153 -7267 -14119 -7233
rect -14081 -7267 -14047 -7233
rect -14009 -7267 -13975 -7233
rect -13937 -7267 -13903 -7233
rect -13865 -7267 -13831 -7233
rect -13793 -7267 -13759 -7233
rect -13721 -7267 -13687 -7233
rect -13649 -7267 -13615 -7233
rect -13577 -7267 -13543 -7233
rect -13505 -7267 -13471 -7233
rect -13433 -7267 -13399 -7233
rect -13361 -7267 -13327 -7233
rect -13289 -7267 -13255 -7233
rect -13217 -7267 -13183 -7233
rect -13145 -7267 -13111 -7233
rect -13073 -7267 -13039 -7233
rect -13001 -7267 -12967 -7233
rect -12929 -7267 -12895 -7233
rect -12857 -7267 -12823 -7233
rect -12785 -7267 -12751 -7233
rect -12713 -7267 -12679 -7233
rect -12641 -7267 -12607 -7233
rect -12569 -7267 -12535 -7233
rect -12497 -7267 -12463 -7233
rect -12425 -7267 -12391 -7233
rect -12353 -7267 -12319 -7233
rect -12281 -7267 -12247 -7233
rect -12209 -7267 -12175 -7233
rect -12137 -7267 -12103 -7233
rect -12065 -7267 -12031 -7233
rect -11993 -7267 -11959 -7233
rect -11921 -7267 -11887 -7233
rect -11849 -7267 -11815 -7233
rect -11777 -7267 -11743 -7233
rect -11705 -7267 -11671 -7233
rect -11633 -7267 -11599 -7233
rect -11561 -7267 -11527 -7233
rect -11489 -7267 -11455 -7233
rect -11417 -7267 -11383 -7233
rect -11345 -7267 -11311 -7233
rect -11273 -7267 -11239 -7233
rect -11201 -7267 -11167 -7233
rect -11129 -7267 -11095 -7233
rect -11057 -7267 -11023 -7233
rect -10985 -7267 -10951 -7233
rect -10913 -7267 -10879 -7233
rect -10841 -7267 -10807 -7233
rect -10769 -7267 -10735 -7233
rect -10697 -7267 -10663 -7233
rect -10625 -7267 -10591 -7233
rect -10553 -7267 -10519 -7233
rect -10481 -7267 -10447 -7233
rect -10409 -7267 -10375 -7233
rect -10337 -7267 -10303 -7233
rect -10265 -7267 -10231 -7233
rect -10193 -7267 -10159 -7233
rect -10121 -7267 -10087 -7233
rect -10049 -7267 -10015 -7233
rect -9977 -7267 -9943 -7233
rect -9905 -7267 -9871 -7233
rect -9833 -7267 -9799 -7233
rect -9761 -7267 -9727 -7233
rect -9689 -7267 -9655 -7233
rect -9617 -7267 -9583 -7233
rect -9545 -7267 -9511 -7233
rect -9473 -7267 -9439 -7233
rect -9401 -7267 -9367 -7233
rect -9329 -7267 -9295 -7233
rect -9257 -7267 -9223 -7233
rect -9185 -7267 -9151 -7233
rect -9113 -7267 -9079 -7233
rect -9041 -7267 -9007 -7233
rect -8969 -7267 -8935 -7233
rect -8897 -7267 -8863 -7233
rect -8825 -7267 -8791 -7233
rect -8753 -7267 -8719 -7233
rect -8681 -7267 -8647 -7233
rect -8609 -7267 -8575 -7233
rect -8537 -7267 -8503 -7233
rect -8465 -7267 -8431 -7233
rect -8393 -7267 -8359 -7233
rect -8321 -7267 -8287 -7233
rect -8249 -7267 -8215 -7233
rect -8177 -7267 -8143 -7233
rect -8105 -7267 -8071 -7233
rect -8033 -7267 -7999 -7233
rect -7961 -7267 -7927 -7233
rect -7889 -7267 -7855 -7233
rect -7817 -7267 -7783 -7233
rect -7745 -7267 -7711 -7233
rect -7673 -7267 -7639 -7233
rect -7601 -7267 -7567 -7233
rect -7529 -7267 -7495 -7233
rect -7457 -7267 -7423 -7233
rect -7385 -7267 -7351 -7233
rect -7313 -7267 -7279 -7233
rect -7241 -7267 -7207 -7233
rect -7169 -7267 -7135 -7233
rect -7097 -7267 -7063 -7233
rect -7025 -7267 -6991 -7233
rect -6953 -7267 -6919 -7233
rect -6881 -7267 -6847 -7233
rect -6809 -7267 -6775 -7233
rect -6737 -7267 -6703 -7233
rect -6665 -7267 -6631 -7233
rect -6593 -7267 -6559 -7233
rect -6521 -7267 -6487 -7233
rect -6449 -7267 -6415 -7233
rect -6377 -7267 -6343 -7233
rect -6305 -7267 -6271 -7233
rect -6233 -7267 -6199 -7233
rect -6161 -7267 -6127 -7233
rect -6089 -7267 -6055 -7233
rect -6017 -7267 -5983 -7233
rect -5945 -7267 -5911 -7233
rect -5873 -7267 -5839 -7233
rect -5801 -7267 -5767 -7233
rect -5729 -7267 -5695 -7233
rect -5657 -7267 -5623 -7233
rect -5585 -7267 -5551 -7233
rect -5513 -7267 -5479 -7233
rect -5441 -7267 -5407 -7233
rect -5369 -7267 -5335 -7233
rect -5297 -7267 -5263 -7233
rect -5225 -7267 -5191 -7233
rect -5153 -7267 -5119 -7233
rect -5081 -7267 -5047 -7233
rect -5009 -7267 -4975 -7233
rect -4937 -7267 -4903 -7233
rect -4865 -7267 -4831 -7233
rect -4793 -7267 -4759 -7233
rect -4721 -7267 -4687 -7233
rect -4649 -7267 -4615 -7233
rect -4577 -7267 -4543 -7233
rect -4505 -7267 -4471 -7233
rect -4433 -7267 -4399 -7233
rect -4361 -7267 -4327 -7233
rect -4289 -7267 -4255 -7233
rect -4217 -7267 -4183 -7233
rect -4145 -7267 -4111 -7233
rect -4073 -7267 -4039 -7233
rect -4001 -7267 -3967 -7233
rect -3929 -7267 -3895 -7233
rect -3857 -7267 -3823 -7233
rect -3785 -7267 -3751 -7233
rect -3713 -7267 -3679 -7233
rect -3641 -7267 -3607 -7233
rect -3569 -7267 -3535 -7233
rect -3497 -7267 -3463 -7233
rect -3425 -7267 -3391 -7233
rect -3353 -7267 -3319 -7233
rect -3281 -7267 -3247 -7233
rect -3209 -7267 -3175 -7233
rect -3137 -7267 -3103 -7233
rect -3065 -7267 -3031 -7233
rect -2993 -7267 -2959 -7233
rect -2921 -7267 -2887 -7233
rect -2849 -7267 -2815 -7233
rect -2777 -7267 -2743 -7233
rect -2705 -7267 -2671 -7233
rect -2633 -7267 -2599 -7233
rect -2561 -7267 -2527 -7233
rect -2489 -7267 -2455 -7233
rect -2417 -7267 -2383 -7233
rect -2345 -7267 -2311 -7233
rect -2273 -7267 -2239 -7233
rect -2201 -7267 -2167 -7233
rect -2129 -7267 -2095 -7233
rect -2057 -7267 -2023 -7233
rect -1985 -7267 -1951 -7233
rect -1913 -7267 -1879 -7233
rect -1841 -7267 -1807 -7233
rect -1769 -7267 -1735 -7233
rect -1697 -7267 -1663 -7233
rect -1625 -7267 -1591 -7233
rect -1553 -7267 -1519 -7233
rect -1481 -7267 -1447 -7233
rect -1409 -7267 -1375 -7233
rect -1337 -7267 -1303 -7233
rect -1265 -7267 -1231 -7233
rect -1193 -7267 -1159 -7233
rect -1121 -7267 -1087 -7233
rect -1049 -7267 -1015 -7233
rect -977 -7267 -943 -7233
rect -905 -7267 -871 -7233
rect -833 -7267 -799 -7233
rect -761 -7267 -727 -7233
rect -689 -7267 -655 -7233
rect -617 -7267 -583 -7233
rect -545 -7267 -511 -7233
rect -473 -7267 -439 -7233
rect -401 -7267 -367 -7233
rect -329 -7267 -295 -7233
rect -257 -7267 -223 -7233
rect -185 -7267 -151 -7233
rect -113 -7267 -79 -7233
rect -41 -7267 -7 -7233
rect 31 -7267 65 -7233
rect 103 -7267 137 -7233
rect 175 -7267 209 -7233
rect 247 -7267 281 -7233
rect 319 -7267 353 -7233
rect 391 -7267 425 -7233
rect 463 -7267 497 -7233
rect 535 -7267 569 -7233
rect 607 -7267 641 -7233
rect 679 -7267 713 -7233
rect 751 -7267 785 -7233
rect 823 -7267 857 -7233
rect 895 -7267 929 -7233
rect 967 -7267 1001 -7233
rect 1039 -7267 1073 -7233
rect 1111 -7267 1145 -7233
rect 1183 -7267 1217 -7233
rect 1255 -7267 1289 -7233
rect 1327 -7267 1361 -7233
rect 1399 -7267 1433 -7233
rect 1471 -7267 1505 -7233
rect 1543 -7267 1577 -7233
rect 1615 -7267 1649 -7233
rect 1687 -7267 1721 -7233
rect 1759 -7267 1793 -7233
rect 1831 -7267 1865 -7233
rect 1903 -7267 1937 -7233
rect 1975 -7267 2009 -7233
rect 2047 -7267 2081 -7233
rect 2119 -7267 2153 -7233
rect 2191 -7267 2225 -7233
rect 2263 -7267 2297 -7233
rect 2335 -7267 2369 -7233
rect 2407 -7267 2441 -7233
rect 2479 -7267 2513 -7233
rect 2551 -7267 2585 -7233
rect 2623 -7267 2657 -7233
rect 2695 -7267 2729 -7233
rect 2767 -7267 2801 -7233
rect 2839 -7267 2873 -7233
rect 2911 -7267 2945 -7233
rect 2983 -7267 3017 -7233
rect 3055 -7267 3089 -7233
rect 3127 -7267 3161 -7233
rect 3199 -7267 3233 -7233
rect 3271 -7267 3305 -7233
rect 3343 -7267 3377 -7233
rect 3415 -7267 3449 -7233
rect 3487 -7267 3521 -7233
rect 3559 -7267 3593 -7233
rect 3631 -7267 3665 -7233
rect 3703 -7267 3737 -7233
rect 3775 -7267 3809 -7233
rect 3847 -7267 3881 -7233
rect 3919 -7267 3953 -7233
rect 3991 -7267 4025 -7233
rect 4063 -7267 4097 -7233
rect 4135 -7267 4169 -7233
rect 4207 -7267 4241 -7233
rect 4279 -7267 4313 -7233
rect 4351 -7267 4385 -7233
rect 4423 -7267 4457 -7233
rect 4495 -7267 4529 -7233
rect 4567 -7267 4601 -7233
rect 4639 -7267 4673 -7233
rect 4711 -7267 4745 -7233
rect 4783 -7267 4817 -7233
rect 4855 -7267 4889 -7233
rect 4927 -7267 4961 -7233
rect 4999 -7267 5033 -7233
rect 5071 -7267 5105 -7233
rect 5143 -7267 5177 -7233
rect 5215 -7267 5249 -7233
rect 5287 -7267 5321 -7233
rect 5359 -7267 5393 -7233
rect 5431 -7267 5465 -7233
rect 5503 -7267 5537 -7233
rect 5575 -7267 5609 -7233
rect 5647 -7267 5681 -7233
rect 5719 -7267 5753 -7233
rect 5791 -7267 5825 -7233
rect 5863 -7267 5897 -7233
rect 5935 -7267 5969 -7233
rect 6007 -7267 6041 -7233
rect 6079 -7267 6113 -7233
rect 6151 -7267 6185 -7233
rect 6223 -7267 6257 -7233
rect 6295 -7267 6329 -7233
rect 6367 -7267 6401 -7233
rect 6439 -7267 6473 -7233
rect 6511 -7267 6545 -7233
rect 6583 -7267 6617 -7233
rect 6655 -7267 6689 -7233
rect 6727 -7267 6761 -7233
rect 6799 -7267 6833 -7233
rect 6871 -7267 6905 -7233
rect 6943 -7267 6977 -7233
rect 7015 -7267 7049 -7233
rect 7087 -7267 7121 -7233
rect 7159 -7267 7193 -7233
rect 7231 -7267 7265 -7233
rect 7303 -7267 7337 -7233
rect 7375 -7267 7409 -7233
rect 7447 -7267 7481 -7233
rect 7519 -7267 7553 -7233
rect 7591 -7267 7625 -7233
rect 7663 -7267 7697 -7233
rect 7735 -7267 7769 -7233
rect 7807 -7267 7841 -7233
rect 7879 -7267 7913 -7233
rect 7951 -7267 7985 -7233
rect 8023 -7267 8057 -7233
rect 8095 -7267 8129 -7233
rect 8167 -7267 8201 -7233
rect 8239 -7267 8273 -7233
rect 8311 -7267 8345 -7233
rect 8383 -7267 8417 -7233
rect 8455 -7267 8489 -7233
rect 8527 -7267 8561 -7233
rect 8599 -7267 8633 -7233
rect 8671 -7267 8705 -7233
rect 8743 -7267 8777 -7233
rect 8815 -7267 8849 -7233
rect 8887 -7267 8921 -7233
rect 8959 -7267 8993 -7233
rect 9031 -7267 9065 -7233
rect 9103 -7267 9137 -7233
rect 9175 -7267 9209 -7233
rect 9247 -7267 9281 -7233
rect 9319 -7267 9353 -7233
rect 9391 -7267 9425 -7233
rect 9463 -7267 9497 -7233
rect 9535 -7267 9569 -7233
rect 9607 -7267 9641 -7233
rect 9679 -7267 9713 -7233
rect 9751 -7267 9785 -7233
rect 9823 -7267 9857 -7233
rect 9895 -7267 9929 -7233
rect 9967 -7267 10001 -7233
rect 10039 -7267 10073 -7233
rect 10111 -7267 10145 -7233
rect 10183 -7267 10217 -7233
rect 10255 -7267 10289 -7233
rect 10327 -7267 10361 -7233
rect 10399 -7267 10433 -7233
rect 10471 -7267 10505 -7233
rect 10543 -7267 10577 -7233
rect 10615 -7267 10649 -7233
rect 10687 -7267 10721 -7233
rect 10759 -7267 10793 -7233
rect 10831 -7267 10865 -7233
rect 10903 -7267 10937 -7233
rect 10975 -7267 11009 -7233
rect 11047 -7267 11081 -7233
rect 11119 -7267 11153 -7233
rect 11191 -7267 11225 -7233
rect 11263 -7267 11297 -7233
rect 11335 -7267 11369 -7233
rect 11407 -7267 11441 -7233
rect 11479 -7267 11513 -7233
rect 11551 -7267 11585 -7233
rect 11623 -7267 11657 -7233
rect 11695 -7267 11729 -7233
rect 11767 -7267 11801 -7233
rect 11839 -7267 11873 -7233
rect 11911 -7267 11945 -7233
rect 11983 -7267 12017 -7233
rect 12055 -7267 12089 -7233
rect 12127 -7267 12161 -7233
rect 12199 -7267 12233 -7233
rect 12271 -7267 12305 -7233
rect 12343 -7267 12377 -7233
rect 12415 -7267 12449 -7233
rect 12487 -7267 12521 -7233
rect 12559 -7267 12593 -7233
rect 12631 -7267 12665 -7233
rect 12703 -7267 12737 -7233
rect 12775 -7267 12809 -7233
rect 12847 -7267 12881 -7233
rect 12919 -7267 12953 -7233
rect 12991 -7267 13025 -7233
rect 13063 -7267 13097 -7233
rect 13135 -7267 13169 -7233
rect 13207 -7267 13241 -7233
rect 13279 -7267 13313 -7233
rect 13351 -7267 13385 -7233
rect 13423 -7267 13457 -7233
rect 13495 -7267 13529 -7233
rect 13567 -7267 13601 -7233
rect 13639 -7267 13673 -7233
rect 13711 -7267 13745 -7233
rect 13783 -7267 13817 -7233
rect 13855 -7267 13889 -7233
rect 13927 -7267 13961 -7233
rect 13999 -7267 14033 -7233
rect 14071 -7267 14105 -7233
rect 14143 -7267 14177 -7233
rect 14215 -7267 14249 -7233
rect 14287 -7267 14321 -7233
rect 14359 -7267 14393 -7233
rect 14431 -7267 14465 -7233
rect 14503 -7267 14537 -7233
rect 14575 -7267 14609 -7233
rect 14647 -7267 14681 -7233
rect 14719 -7267 14753 -7233
rect 14791 -7267 14825 -7233
rect 14863 -7267 14897 -7233
rect 14935 -7267 14969 -7233
rect 15007 -7267 15041 -7233
rect 15079 -7267 15113 -7233
rect 15151 -7267 15185 -7233
rect 15223 -7267 15257 -7233
rect 15295 -7267 15329 -7233
rect 15367 -7267 15401 -7233
rect 15439 -7267 15473 -7233
rect 15511 -7267 15545 -7233
rect 15583 -7267 15617 -7233
rect 15655 -7267 15689 -7233
rect 15727 -7267 15761 -7233
rect 15799 -7267 15833 -7233
rect 15871 -7267 15905 -7233
rect 15943 -7267 15977 -7233
rect 16015 -7267 16049 -7233
rect 16087 -7267 16121 -7233
rect 16159 -7267 16193 -7233
rect 16231 -7267 16265 -7233
rect 16303 -7267 16337 -7233
rect 16375 -7267 16409 -7233
rect 16447 -7267 16481 -7233
rect 16519 -7267 16553 -7233
rect 16591 -7267 16625 -7233
rect 16663 -7267 16697 -7233
rect 16735 -7267 16769 -7233
rect 16807 -7267 16841 -7233
rect 16879 -7267 16913 -7233
rect 16951 -7267 16985 -7233
rect 17023 -7267 17057 -7233
rect 17095 -7267 17129 -7233
rect 17167 -7267 17201 -7233
rect 17239 -7267 17273 -7233
rect 17311 -7267 17345 -7233
rect 17383 -7267 17417 -7233
rect 17455 -7267 17489 -7233
rect 17527 -7267 17561 -7233
rect 17599 -7267 17633 -7233
rect 17671 -7267 17705 -7233
rect 17743 -7267 17777 -7233
rect 17815 -7267 17849 -7233
rect 17887 -7267 17921 -7233
rect 17959 -7267 17993 -7233
rect 18031 -7267 18065 -7233
rect 18103 -7267 18137 -7233
rect 18175 -7267 18209 -7233
rect 18247 -7267 18281 -7233
rect 18319 -7267 18353 -7233
rect 18391 -7267 18425 -7233
rect 18463 -7267 18497 -7233
rect 18535 -7267 18569 -7233
rect 18607 -7267 18641 -7233
rect 18679 -7267 18713 -7233
rect 18751 -7267 18785 -7233
rect 18823 -7267 18857 -7233
rect 18895 -7267 18929 -7233
rect 18967 -7267 19001 -7233
rect 19039 -7267 19073 -7233
rect 19111 -7267 19145 -7233
rect 19183 -7267 19217 -7233
rect 19255 -7267 19289 -7233
rect 19327 -7267 19361 -7233
rect 19399 -7267 19433 -7233
rect 19471 -7267 19505 -7233
rect 19543 -7267 19577 -7233
rect 19615 -7267 19649 -7233
rect 19687 -7267 19721 -7233
rect 19759 -7267 19793 -7233
rect 19831 -7267 19865 -7233
rect 19903 -7267 19937 -7233
rect 19975 -7267 20009 -7233
rect 20047 -7267 20081 -7233
rect 20119 -7267 20153 -7233
rect 20191 -7267 20225 -7233
rect 20263 -7267 20297 -7233
rect 20335 -7267 20369 -7233
rect 20407 -7267 20441 -7233
rect 20479 -7267 20513 -7233
rect 20551 -7267 20585 -7233
rect 20623 -7267 20657 -7233
rect 20695 -7267 20729 -7233
rect 20767 -7267 20801 -7233
rect 20839 -7267 20873 -7233
rect 20911 -7267 20945 -7233
rect 20983 -7267 21017 -7233
rect 21055 -7267 21089 -7233
rect 21127 -7267 21161 -7233
rect 21199 -7267 21233 -7233
rect 21271 -7267 21305 -7233
rect 21343 -7267 21377 -7233
rect 21415 -7267 21449 -7233
rect 21487 -7267 21521 -7233
rect 21559 -7267 21593 -7233
rect 21631 -7267 21665 -7233
rect 21703 -7267 21737 -7233
rect 21775 -7267 21809 -7233
rect 21847 -7267 21881 -7233
rect 21919 -7267 21953 -7233
rect 21991 -7267 22025 -7233
rect 22063 -7267 22097 -7233
rect 22135 -7267 22169 -7233
rect 22207 -7267 22241 -7233
rect 22279 -7267 22313 -7233
rect 22351 -7267 22385 -7233
rect 22423 -7267 22457 -7233
rect 22495 -7267 22529 -7233
rect 22567 -7267 22601 -7233
rect 22639 -7267 22673 -7233
rect 22711 -7267 22745 -7233
rect 22783 -7267 22817 -7233
rect 22855 -7267 22889 -7233
rect 22927 -7267 22961 -7233
rect 22999 -7267 23033 -7233
rect 23071 -7267 23105 -7233
rect 23143 -7267 23177 -7233
rect 23215 -7267 23249 -7233
rect 23287 -7267 23321 -7233
rect 23359 -7267 23393 -7233
rect 23431 -7267 23465 -7233
rect 23503 -7267 23537 -7233
rect 23575 -7267 23609 -7233
rect 23647 -7267 23681 -7233
rect 23719 -7267 23753 -7233
rect 23791 -7267 23825 -7233
rect 23863 -7267 23897 -7233
rect 23935 -7267 23969 -7233
rect 24007 -7267 24041 -7233
rect 24079 -7267 24113 -7233
rect 24151 -7267 24185 -7233
rect 24223 -7267 24257 -7233
rect 24295 -7267 24329 -7233
rect 24367 -7267 24401 -7233
rect 24439 -7267 24473 -7233
rect 24511 -7267 24545 -7233
rect 24583 -7267 24617 -7233
rect 24655 -7267 24689 -7233
rect 24727 -7267 24761 -7233
rect 24799 -7267 24833 -7233
rect 24871 -7267 24905 -7233
rect 24943 -7267 24977 -7233
rect 25015 -7267 25049 -7233
rect 25087 -7267 25121 -7233
rect 25159 -7267 25193 -7233
rect 25231 -7267 25265 -7233
rect 25303 -7267 25337 -7233
rect 25375 -7267 25409 -7233
rect 25447 -7267 25481 -7233
rect 25519 -7267 25553 -7233
rect 25591 -7267 25625 -7233
rect 25663 -7267 25697 -7233
rect 25735 -7267 25769 -7233
rect 25807 -7267 25841 -7233
rect 25879 -7267 25913 -7233
rect 25951 -7267 25985 -7233
rect 26023 -7267 26057 -7233
rect 26095 -7267 26129 -7233
rect 26167 -7267 26201 -7233
rect 26239 -7267 26273 -7233
rect 26311 -7267 26345 -7233
rect 26383 -7267 26417 -7233
rect 26455 -7267 26489 -7233
rect 26527 -7267 26561 -7233
rect 26599 -7267 26633 -7233
rect 26671 -7267 26705 -7233
rect 26743 -7267 26777 -7233
rect 26815 -7267 26849 -7233
rect 26887 -7267 26921 -7233
rect 26959 -7267 26993 -7233
rect 27031 -7267 27065 -7233
rect 27103 -7267 27137 -7233
rect 27175 -7267 27209 -7233
rect 27247 -7267 27281 -7233
rect 27319 -7267 27353 -7233
rect 27391 -7267 27425 -7233
rect 27463 -7267 27497 -7233
rect 27535 -7267 27569 -7233
rect 27607 -7267 27641 -7233
rect 27679 -7267 27713 -7233
rect 27751 -7267 27785 -7233
rect 27823 -7267 27857 -7233
rect 27895 -7267 27929 -7233
rect 27967 -7267 28001 -7233
rect 28039 -7267 28073 -7233
rect 28111 -7267 28145 -7233
rect 28183 -7267 28217 -7233
rect 28255 -7267 28289 -7233
rect 28327 -7267 28361 -7233
rect 28399 -7267 28433 -7233
rect 28471 -7267 28505 -7233
rect 28543 -7267 28577 -7233
rect 28615 -7267 28649 -7233
rect 28687 -7267 28721 -7233
rect 28759 -7267 28793 -7233
rect 28831 -7267 28865 -7233
rect 28903 -7267 28937 -7233
rect 28975 -7267 29009 -7233
rect 29047 -7267 29081 -7233
rect 29119 -7267 29153 -7233
rect 29191 -7267 29225 -7233
rect 29263 -7267 29297 -7233
rect 29335 -7267 29369 -7233
rect 29407 -7267 29441 -7233
rect 29479 -7267 29513 -7233
rect 29551 -7267 29585 -7233
rect 29623 -7267 29657 -7233
rect 29695 -7267 29729 -7233
rect 29767 -7267 29801 -7233
rect 29839 -7267 29873 -7233
rect 29911 -7267 29945 -7233
rect 29983 -7267 30017 -7233
rect 30055 -7267 30089 -7233
rect 30127 -7267 30161 -7233
rect 30199 -7267 30233 -7233
rect 30271 -7267 30305 -7233
rect 30343 -7267 30377 -7233
rect 30415 -7267 30449 -7233
rect 30487 -7267 30521 -7233
rect 30559 -7267 30593 -7233
rect 30631 -7267 30665 -7233
rect 30703 -7267 30737 -7233
rect 30775 -7267 30809 -7233
rect 30847 -7267 30881 -7233
rect 30919 -7267 30953 -7233
rect 30991 -7267 31025 -7233
rect 31063 -7267 31097 -7233
rect 31135 -7267 31169 -7233
rect 31207 -7267 31241 -7233
rect 31279 -7267 31313 -7233
rect 31351 -7267 31385 -7233
rect 31423 -7267 31457 -7233
rect 31495 -7267 31529 -7233
rect 31567 -7267 31601 -7233
rect 31639 -7267 31673 -7233
rect 31711 -7267 31745 -7233
rect 31783 -7267 31817 -7233
rect 31855 -7267 31889 -7233
rect 31927 -7267 31961 -7233
rect 31999 -7267 32033 -7233
rect 32071 -7267 32105 -7233
rect 32143 -7267 32177 -7233
rect 32215 -7267 32249 -7233
rect 32287 -7267 32321 -7233
rect 32359 -7267 32393 -7233
rect 32431 -7267 32465 -7233
rect 32503 -7267 32537 -7233
rect 32575 -7267 32609 -7233
rect 32647 -7267 32681 -7233
rect 32719 -7267 32753 -7233
rect 32791 -7267 32825 -7233
rect 32863 -7267 32897 -7233
rect 32935 -7267 32969 -7233
rect 33007 -7267 33041 -7233
rect 33079 -7267 33113 -7233
rect 33151 -7267 33185 -7233
rect 33223 -7267 33257 -7233
rect 33295 -7267 33329 -7233
rect 33367 -7267 33401 -7233
rect 33439 -7267 33473 -7233
rect 33511 -7267 33545 -7233
rect 33583 -7267 33617 -7233
rect 33655 -7267 33689 -7233
rect 33727 -7267 33761 -7233
rect 33799 -7267 33833 -7233
rect 33871 -7267 33905 -7233
rect 33943 -7267 33977 -7233
rect 34015 -7267 34049 -7233
rect 34087 -7267 34121 -7233
rect 34159 -7267 34193 -7233
rect 34231 -7267 34265 -7233
rect 34303 -7267 34337 -7233
rect 34375 -7267 34409 -7233
rect 34447 -7267 34481 -7233
rect 34519 -7267 34553 -7233
rect 34591 -7267 34625 -7233
rect 34663 -7267 34697 -7233
rect 34735 -7267 34769 -7233
rect 34807 -7267 34841 -7233
rect 34879 -7267 34913 -7233
rect 34951 -7267 34985 -7233
rect 35023 -7267 35057 -7233
rect 35095 -7267 35129 -7233
rect 35167 -7267 35201 -7233
<< metal1 >>
rect -17500 14867 35400 14900
rect -17500 14833 -17301 14867
rect -17267 14833 -17229 14867
rect -17195 14833 -17157 14867
rect -17123 14833 -17085 14867
rect -17051 14833 -17013 14867
rect -16979 14833 -16941 14867
rect -16907 14833 -16869 14867
rect -16835 14833 -16797 14867
rect -16763 14833 -16725 14867
rect -16691 14833 -16653 14867
rect -16619 14833 -16581 14867
rect -16547 14833 -16509 14867
rect -16475 14833 -16437 14867
rect -16403 14833 -16365 14867
rect -16331 14833 -16293 14867
rect -16259 14833 -16221 14867
rect -16187 14833 -16149 14867
rect -16115 14833 -16077 14867
rect -16043 14833 -16005 14867
rect -15971 14833 -15933 14867
rect -15899 14833 -15861 14867
rect -15827 14833 -15789 14867
rect -15755 14833 -15717 14867
rect -15683 14833 -15645 14867
rect -15611 14833 -15573 14867
rect -15539 14833 -15501 14867
rect -15467 14833 -15429 14867
rect -15395 14833 -15357 14867
rect -15323 14833 -15285 14867
rect -15251 14833 -15213 14867
rect -15179 14833 -15141 14867
rect -15107 14833 -15069 14867
rect -15035 14833 -14997 14867
rect -14963 14833 -14925 14867
rect -14891 14833 -14853 14867
rect -14819 14833 -14781 14867
rect -14747 14833 -14709 14867
rect -14675 14833 -14637 14867
rect -14603 14833 -14565 14867
rect -14531 14833 -14493 14867
rect -14459 14833 -14421 14867
rect -14387 14833 -14349 14867
rect -14315 14833 -14277 14867
rect -14243 14833 -14205 14867
rect -14171 14833 -14133 14867
rect -14099 14833 -14061 14867
rect -14027 14833 -13989 14867
rect -13955 14833 -13917 14867
rect -13883 14833 -13845 14867
rect -13811 14833 -13773 14867
rect -13739 14833 -13701 14867
rect -13667 14833 -13629 14867
rect -13595 14833 -13557 14867
rect -13523 14833 -13485 14867
rect -13451 14833 -13413 14867
rect -13379 14833 -13341 14867
rect -13307 14833 -13269 14867
rect -13235 14833 -13197 14867
rect -13163 14833 -13125 14867
rect -13091 14833 -13053 14867
rect -13019 14833 -12981 14867
rect -12947 14833 -12909 14867
rect -12875 14833 -12837 14867
rect -12803 14833 -12765 14867
rect -12731 14833 -12693 14867
rect -12659 14833 -12621 14867
rect -12587 14833 -12549 14867
rect -12515 14833 -12477 14867
rect -12443 14833 -12405 14867
rect -12371 14833 -12333 14867
rect -12299 14833 -12261 14867
rect -12227 14833 -12189 14867
rect -12155 14833 -12117 14867
rect -12083 14833 -12045 14867
rect -12011 14833 -11973 14867
rect -11939 14833 -11901 14867
rect -11867 14833 -11829 14867
rect -11795 14833 -11757 14867
rect -11723 14833 -11685 14867
rect -11651 14833 -11613 14867
rect -11579 14833 -11541 14867
rect -11507 14833 -11469 14867
rect -11435 14833 -11397 14867
rect -11363 14833 -11325 14867
rect -11291 14833 -11253 14867
rect -11219 14833 -11181 14867
rect -11147 14833 -11109 14867
rect -11075 14833 -11037 14867
rect -11003 14833 -10965 14867
rect -10931 14833 -10893 14867
rect -10859 14833 -10821 14867
rect -10787 14833 -10749 14867
rect -10715 14833 -10677 14867
rect -10643 14833 -10605 14867
rect -10571 14833 -10533 14867
rect -10499 14833 -10461 14867
rect -10427 14833 -10389 14867
rect -10355 14833 -10317 14867
rect -10283 14833 -10245 14867
rect -10211 14833 -10173 14867
rect -10139 14833 -10101 14867
rect -10067 14833 -10029 14867
rect -9995 14833 -9957 14867
rect -9923 14833 -9885 14867
rect -9851 14833 -9813 14867
rect -9779 14833 -9741 14867
rect -9707 14833 -9669 14867
rect -9635 14833 -9597 14867
rect -9563 14833 -9525 14867
rect -9491 14833 -9453 14867
rect -9419 14833 -9381 14867
rect -9347 14833 -9309 14867
rect -9275 14833 -9237 14867
rect -9203 14833 -9165 14867
rect -9131 14833 -9093 14867
rect -9059 14833 -9021 14867
rect -8987 14833 -8949 14867
rect -8915 14833 -8877 14867
rect -8843 14833 -8805 14867
rect -8771 14833 -8733 14867
rect -8699 14833 -8661 14867
rect -8627 14833 -8589 14867
rect -8555 14833 -8517 14867
rect -8483 14833 -8445 14867
rect -8411 14833 -8373 14867
rect -8339 14833 -8301 14867
rect -8267 14833 -8229 14867
rect -8195 14833 -8157 14867
rect -8123 14833 -8085 14867
rect -8051 14833 -8013 14867
rect -7979 14833 -7941 14867
rect -7907 14833 -7869 14867
rect -7835 14833 -7797 14867
rect -7763 14833 -7725 14867
rect -7691 14833 -7653 14867
rect -7619 14833 -7581 14867
rect -7547 14833 -7509 14867
rect -7475 14833 -7437 14867
rect -7403 14833 -7365 14867
rect -7331 14833 -7293 14867
rect -7259 14833 -7221 14867
rect -7187 14833 -7149 14867
rect -7115 14833 -7077 14867
rect -7043 14833 -7005 14867
rect -6971 14833 -6933 14867
rect -6899 14833 -6861 14867
rect -6827 14833 -6789 14867
rect -6755 14833 -6717 14867
rect -6683 14833 -6645 14867
rect -6611 14833 -6573 14867
rect -6539 14833 -6501 14867
rect -6467 14833 -6429 14867
rect -6395 14833 -6357 14867
rect -6323 14833 -6285 14867
rect -6251 14833 -6213 14867
rect -6179 14833 -6141 14867
rect -6107 14833 -6069 14867
rect -6035 14833 -5997 14867
rect -5963 14833 -5925 14867
rect -5891 14833 -5853 14867
rect -5819 14833 -5781 14867
rect -5747 14833 -5709 14867
rect -5675 14833 -5637 14867
rect -5603 14833 -5565 14867
rect -5531 14833 -5493 14867
rect -5459 14833 -5421 14867
rect -5387 14833 -5349 14867
rect -5315 14833 -5277 14867
rect -5243 14833 -5205 14867
rect -5171 14833 -5133 14867
rect -5099 14833 -5061 14867
rect -5027 14833 -4989 14867
rect -4955 14833 -4917 14867
rect -4883 14833 -4845 14867
rect -4811 14833 -4773 14867
rect -4739 14833 -4701 14867
rect -4667 14833 -4629 14867
rect -4595 14833 -4557 14867
rect -4523 14833 -4485 14867
rect -4451 14833 -4413 14867
rect -4379 14833 -4341 14867
rect -4307 14833 -4269 14867
rect -4235 14833 -4197 14867
rect -4163 14833 -4125 14867
rect -4091 14833 -4053 14867
rect -4019 14833 -3981 14867
rect -3947 14833 -3909 14867
rect -3875 14833 -3837 14867
rect -3803 14833 -3765 14867
rect -3731 14833 -3693 14867
rect -3659 14833 -3621 14867
rect -3587 14833 -3549 14867
rect -3515 14833 -3477 14867
rect -3443 14833 -3405 14867
rect -3371 14833 -3333 14867
rect -3299 14833 -3261 14867
rect -3227 14833 -3189 14867
rect -3155 14833 -3117 14867
rect -3083 14833 -3045 14867
rect -3011 14833 -2973 14867
rect -2939 14833 -2901 14867
rect -2867 14833 -2829 14867
rect -2795 14833 -2757 14867
rect -2723 14833 -2685 14867
rect -2651 14833 -2613 14867
rect -2579 14833 -2541 14867
rect -2507 14833 -2469 14867
rect -2435 14833 -2397 14867
rect -2363 14833 -2325 14867
rect -2291 14833 -2253 14867
rect -2219 14833 -2181 14867
rect -2147 14833 -2109 14867
rect -2075 14833 -2037 14867
rect -2003 14833 -1965 14867
rect -1931 14833 -1893 14867
rect -1859 14833 -1821 14867
rect -1787 14833 -1749 14867
rect -1715 14833 -1677 14867
rect -1643 14833 -1605 14867
rect -1571 14833 -1533 14867
rect -1499 14833 -1461 14867
rect -1427 14833 -1389 14867
rect -1355 14833 -1317 14867
rect -1283 14833 -1245 14867
rect -1211 14833 -1173 14867
rect -1139 14833 -1101 14867
rect -1067 14833 -1029 14867
rect -995 14833 -957 14867
rect -923 14833 -885 14867
rect -851 14833 -813 14867
rect -779 14833 -741 14867
rect -707 14833 -669 14867
rect -635 14833 -597 14867
rect -563 14833 -525 14867
rect -491 14833 -453 14867
rect -419 14833 -381 14867
rect -347 14833 -309 14867
rect -275 14833 -237 14867
rect -203 14833 -165 14867
rect -131 14833 -93 14867
rect -59 14833 -21 14867
rect 13 14833 51 14867
rect 85 14833 123 14867
rect 157 14833 195 14867
rect 229 14833 267 14867
rect 301 14833 339 14867
rect 373 14833 411 14867
rect 445 14833 483 14867
rect 517 14833 555 14867
rect 589 14833 627 14867
rect 661 14833 699 14867
rect 733 14833 771 14867
rect 805 14833 843 14867
rect 877 14833 915 14867
rect 949 14833 987 14867
rect 1021 14833 1059 14867
rect 1093 14833 1131 14867
rect 1165 14833 1203 14867
rect 1237 14833 1275 14867
rect 1309 14833 1347 14867
rect 1381 14833 1419 14867
rect 1453 14833 1491 14867
rect 1525 14833 1563 14867
rect 1597 14833 1635 14867
rect 1669 14833 1707 14867
rect 1741 14833 1779 14867
rect 1813 14833 1851 14867
rect 1885 14833 1923 14867
rect 1957 14833 1995 14867
rect 2029 14833 2067 14867
rect 2101 14833 2139 14867
rect 2173 14833 2211 14867
rect 2245 14833 2283 14867
rect 2317 14833 2355 14867
rect 2389 14833 2427 14867
rect 2461 14833 2499 14867
rect 2533 14833 2571 14867
rect 2605 14833 2643 14867
rect 2677 14833 2715 14867
rect 2749 14833 2787 14867
rect 2821 14833 2859 14867
rect 2893 14833 2931 14867
rect 2965 14833 3003 14867
rect 3037 14833 3075 14867
rect 3109 14833 3147 14867
rect 3181 14833 3219 14867
rect 3253 14833 3291 14867
rect 3325 14833 3363 14867
rect 3397 14833 3435 14867
rect 3469 14833 3507 14867
rect 3541 14833 3579 14867
rect 3613 14833 3651 14867
rect 3685 14833 3723 14867
rect 3757 14833 3795 14867
rect 3829 14833 3867 14867
rect 3901 14833 3939 14867
rect 3973 14833 4011 14867
rect 4045 14833 4083 14867
rect 4117 14833 4155 14867
rect 4189 14833 4227 14867
rect 4261 14833 4299 14867
rect 4333 14833 4371 14867
rect 4405 14833 4443 14867
rect 4477 14833 4515 14867
rect 4549 14833 4587 14867
rect 4621 14833 4659 14867
rect 4693 14833 4731 14867
rect 4765 14833 4803 14867
rect 4837 14833 4875 14867
rect 4909 14833 4947 14867
rect 4981 14833 5019 14867
rect 5053 14833 5091 14867
rect 5125 14833 5163 14867
rect 5197 14833 5235 14867
rect 5269 14833 5307 14867
rect 5341 14833 5379 14867
rect 5413 14833 5451 14867
rect 5485 14833 5523 14867
rect 5557 14833 5595 14867
rect 5629 14833 5667 14867
rect 5701 14833 5739 14867
rect 5773 14833 5811 14867
rect 5845 14833 5883 14867
rect 5917 14833 5955 14867
rect 5989 14833 6027 14867
rect 6061 14833 6099 14867
rect 6133 14833 6171 14867
rect 6205 14833 6243 14867
rect 6277 14833 6315 14867
rect 6349 14833 6387 14867
rect 6421 14833 6459 14867
rect 6493 14833 6531 14867
rect 6565 14833 6603 14867
rect 6637 14833 6675 14867
rect 6709 14833 6747 14867
rect 6781 14833 6819 14867
rect 6853 14833 6891 14867
rect 6925 14833 6963 14867
rect 6997 14833 7035 14867
rect 7069 14833 7107 14867
rect 7141 14833 7179 14867
rect 7213 14833 7251 14867
rect 7285 14833 7323 14867
rect 7357 14833 7395 14867
rect 7429 14833 7467 14867
rect 7501 14833 7539 14867
rect 7573 14833 7611 14867
rect 7645 14833 7683 14867
rect 7717 14833 7755 14867
rect 7789 14833 7827 14867
rect 7861 14833 7899 14867
rect 7933 14833 7971 14867
rect 8005 14833 8043 14867
rect 8077 14833 8115 14867
rect 8149 14833 8187 14867
rect 8221 14833 8259 14867
rect 8293 14833 8331 14867
rect 8365 14833 8403 14867
rect 8437 14833 8475 14867
rect 8509 14833 8547 14867
rect 8581 14833 8619 14867
rect 8653 14833 8691 14867
rect 8725 14833 8763 14867
rect 8797 14833 8835 14867
rect 8869 14833 8907 14867
rect 8941 14833 8979 14867
rect 9013 14833 9051 14867
rect 9085 14833 9123 14867
rect 9157 14833 9195 14867
rect 9229 14833 9267 14867
rect 9301 14833 9339 14867
rect 9373 14833 9411 14867
rect 9445 14833 9483 14867
rect 9517 14833 9555 14867
rect 9589 14833 9627 14867
rect 9661 14833 9699 14867
rect 9733 14833 9771 14867
rect 9805 14833 9843 14867
rect 9877 14833 9915 14867
rect 9949 14833 9987 14867
rect 10021 14833 10059 14867
rect 10093 14833 10131 14867
rect 10165 14833 10203 14867
rect 10237 14833 10275 14867
rect 10309 14833 10347 14867
rect 10381 14833 10419 14867
rect 10453 14833 10491 14867
rect 10525 14833 10563 14867
rect 10597 14833 10635 14867
rect 10669 14833 10707 14867
rect 10741 14833 10779 14867
rect 10813 14833 10851 14867
rect 10885 14833 10923 14867
rect 10957 14833 10995 14867
rect 11029 14833 11067 14867
rect 11101 14833 11139 14867
rect 11173 14833 11211 14867
rect 11245 14833 11283 14867
rect 11317 14833 11355 14867
rect 11389 14833 11427 14867
rect 11461 14833 11499 14867
rect 11533 14833 11571 14867
rect 11605 14833 11643 14867
rect 11677 14833 11715 14867
rect 11749 14833 11787 14867
rect 11821 14833 11859 14867
rect 11893 14833 11931 14867
rect 11965 14833 12003 14867
rect 12037 14833 12075 14867
rect 12109 14833 12147 14867
rect 12181 14833 12219 14867
rect 12253 14833 12291 14867
rect 12325 14833 12363 14867
rect 12397 14833 12435 14867
rect 12469 14833 12507 14867
rect 12541 14833 12579 14867
rect 12613 14833 12651 14867
rect 12685 14833 12723 14867
rect 12757 14833 12795 14867
rect 12829 14833 12867 14867
rect 12901 14833 12939 14867
rect 12973 14833 13011 14867
rect 13045 14833 13083 14867
rect 13117 14833 13155 14867
rect 13189 14833 13227 14867
rect 13261 14833 13299 14867
rect 13333 14833 13371 14867
rect 13405 14833 13443 14867
rect 13477 14833 13515 14867
rect 13549 14833 13587 14867
rect 13621 14833 13659 14867
rect 13693 14833 13731 14867
rect 13765 14833 13803 14867
rect 13837 14833 13875 14867
rect 13909 14833 13947 14867
rect 13981 14833 14019 14867
rect 14053 14833 14091 14867
rect 14125 14833 14163 14867
rect 14197 14833 14235 14867
rect 14269 14833 14307 14867
rect 14341 14833 14379 14867
rect 14413 14833 14451 14867
rect 14485 14833 14523 14867
rect 14557 14833 14595 14867
rect 14629 14833 14667 14867
rect 14701 14833 14739 14867
rect 14773 14833 14811 14867
rect 14845 14833 14883 14867
rect 14917 14833 14955 14867
rect 14989 14833 15027 14867
rect 15061 14833 15099 14867
rect 15133 14833 15171 14867
rect 15205 14833 15243 14867
rect 15277 14833 15315 14867
rect 15349 14833 15387 14867
rect 15421 14833 15459 14867
rect 15493 14833 15531 14867
rect 15565 14833 15603 14867
rect 15637 14833 15675 14867
rect 15709 14833 15747 14867
rect 15781 14833 15819 14867
rect 15853 14833 15891 14867
rect 15925 14833 15963 14867
rect 15997 14833 16035 14867
rect 16069 14833 16107 14867
rect 16141 14833 16179 14867
rect 16213 14833 16251 14867
rect 16285 14833 16323 14867
rect 16357 14833 16395 14867
rect 16429 14833 16467 14867
rect 16501 14833 16539 14867
rect 16573 14833 16611 14867
rect 16645 14833 16683 14867
rect 16717 14833 16755 14867
rect 16789 14833 16827 14867
rect 16861 14833 16899 14867
rect 16933 14833 16971 14867
rect 17005 14833 17043 14867
rect 17077 14833 17115 14867
rect 17149 14833 17187 14867
rect 17221 14833 17259 14867
rect 17293 14833 17331 14867
rect 17365 14833 17403 14867
rect 17437 14833 17475 14867
rect 17509 14833 17547 14867
rect 17581 14833 17619 14867
rect 17653 14833 17691 14867
rect 17725 14833 17763 14867
rect 17797 14833 17835 14867
rect 17869 14833 17907 14867
rect 17941 14833 17979 14867
rect 18013 14833 18051 14867
rect 18085 14833 18123 14867
rect 18157 14833 18195 14867
rect 18229 14833 18267 14867
rect 18301 14833 18339 14867
rect 18373 14833 18411 14867
rect 18445 14833 18483 14867
rect 18517 14833 18555 14867
rect 18589 14833 18627 14867
rect 18661 14833 18699 14867
rect 18733 14833 18771 14867
rect 18805 14833 18843 14867
rect 18877 14833 18915 14867
rect 18949 14833 18987 14867
rect 19021 14833 19059 14867
rect 19093 14833 19131 14867
rect 19165 14833 19203 14867
rect 19237 14833 19275 14867
rect 19309 14833 19347 14867
rect 19381 14833 19419 14867
rect 19453 14833 19491 14867
rect 19525 14833 19563 14867
rect 19597 14833 19635 14867
rect 19669 14833 19707 14867
rect 19741 14833 19779 14867
rect 19813 14833 19851 14867
rect 19885 14833 19923 14867
rect 19957 14833 19995 14867
rect 20029 14833 20067 14867
rect 20101 14833 20139 14867
rect 20173 14833 20211 14867
rect 20245 14833 20283 14867
rect 20317 14833 20355 14867
rect 20389 14833 20427 14867
rect 20461 14833 20499 14867
rect 20533 14833 20571 14867
rect 20605 14833 20643 14867
rect 20677 14833 20715 14867
rect 20749 14833 20787 14867
rect 20821 14833 20859 14867
rect 20893 14833 20931 14867
rect 20965 14833 21003 14867
rect 21037 14833 21075 14867
rect 21109 14833 21147 14867
rect 21181 14833 21219 14867
rect 21253 14833 21291 14867
rect 21325 14833 21363 14867
rect 21397 14833 21435 14867
rect 21469 14833 21507 14867
rect 21541 14833 21579 14867
rect 21613 14833 21651 14867
rect 21685 14833 21723 14867
rect 21757 14833 21795 14867
rect 21829 14833 21867 14867
rect 21901 14833 21939 14867
rect 21973 14833 22011 14867
rect 22045 14833 22083 14867
rect 22117 14833 22155 14867
rect 22189 14833 22227 14867
rect 22261 14833 22299 14867
rect 22333 14833 22371 14867
rect 22405 14833 22443 14867
rect 22477 14833 22515 14867
rect 22549 14833 22587 14867
rect 22621 14833 22659 14867
rect 22693 14833 22731 14867
rect 22765 14833 22803 14867
rect 22837 14833 22875 14867
rect 22909 14833 22947 14867
rect 22981 14833 23019 14867
rect 23053 14833 23091 14867
rect 23125 14833 23163 14867
rect 23197 14833 23235 14867
rect 23269 14833 23307 14867
rect 23341 14833 23379 14867
rect 23413 14833 23451 14867
rect 23485 14833 23523 14867
rect 23557 14833 23595 14867
rect 23629 14833 23667 14867
rect 23701 14833 23739 14867
rect 23773 14833 23811 14867
rect 23845 14833 23883 14867
rect 23917 14833 23955 14867
rect 23989 14833 24027 14867
rect 24061 14833 24099 14867
rect 24133 14833 24171 14867
rect 24205 14833 24243 14867
rect 24277 14833 24315 14867
rect 24349 14833 24387 14867
rect 24421 14833 24459 14867
rect 24493 14833 24531 14867
rect 24565 14833 24603 14867
rect 24637 14833 24675 14867
rect 24709 14833 24747 14867
rect 24781 14833 24819 14867
rect 24853 14833 24891 14867
rect 24925 14833 24963 14867
rect 24997 14833 25035 14867
rect 25069 14833 25107 14867
rect 25141 14833 25179 14867
rect 25213 14833 25251 14867
rect 25285 14833 25323 14867
rect 25357 14833 25395 14867
rect 25429 14833 25467 14867
rect 25501 14833 25539 14867
rect 25573 14833 25611 14867
rect 25645 14833 25683 14867
rect 25717 14833 25755 14867
rect 25789 14833 25827 14867
rect 25861 14833 25899 14867
rect 25933 14833 25971 14867
rect 26005 14833 26043 14867
rect 26077 14833 26115 14867
rect 26149 14833 26187 14867
rect 26221 14833 26259 14867
rect 26293 14833 26331 14867
rect 26365 14833 26403 14867
rect 26437 14833 26475 14867
rect 26509 14833 26547 14867
rect 26581 14833 26619 14867
rect 26653 14833 26691 14867
rect 26725 14833 26763 14867
rect 26797 14833 26835 14867
rect 26869 14833 26907 14867
rect 26941 14833 26979 14867
rect 27013 14833 27051 14867
rect 27085 14833 27123 14867
rect 27157 14833 27195 14867
rect 27229 14833 27267 14867
rect 27301 14833 27339 14867
rect 27373 14833 27411 14867
rect 27445 14833 27483 14867
rect 27517 14833 27555 14867
rect 27589 14833 27627 14867
rect 27661 14833 27699 14867
rect 27733 14833 27771 14867
rect 27805 14833 27843 14867
rect 27877 14833 27915 14867
rect 27949 14833 27987 14867
rect 28021 14833 28059 14867
rect 28093 14833 28131 14867
rect 28165 14833 28203 14867
rect 28237 14833 28275 14867
rect 28309 14833 28347 14867
rect 28381 14833 28419 14867
rect 28453 14833 28491 14867
rect 28525 14833 28563 14867
rect 28597 14833 28635 14867
rect 28669 14833 28707 14867
rect 28741 14833 28779 14867
rect 28813 14833 28851 14867
rect 28885 14833 28923 14867
rect 28957 14833 28995 14867
rect 29029 14833 29067 14867
rect 29101 14833 29139 14867
rect 29173 14833 29211 14867
rect 29245 14833 29283 14867
rect 29317 14833 29355 14867
rect 29389 14833 29427 14867
rect 29461 14833 29499 14867
rect 29533 14833 29571 14867
rect 29605 14833 29643 14867
rect 29677 14833 29715 14867
rect 29749 14833 29787 14867
rect 29821 14833 29859 14867
rect 29893 14833 29931 14867
rect 29965 14833 30003 14867
rect 30037 14833 30075 14867
rect 30109 14833 30147 14867
rect 30181 14833 30219 14867
rect 30253 14833 30291 14867
rect 30325 14833 30363 14867
rect 30397 14833 30435 14867
rect 30469 14833 30507 14867
rect 30541 14833 30579 14867
rect 30613 14833 30651 14867
rect 30685 14833 30723 14867
rect 30757 14833 30795 14867
rect 30829 14833 30867 14867
rect 30901 14833 30939 14867
rect 30973 14833 31011 14867
rect 31045 14833 31083 14867
rect 31117 14833 31155 14867
rect 31189 14833 31227 14867
rect 31261 14833 31299 14867
rect 31333 14833 31371 14867
rect 31405 14833 31443 14867
rect 31477 14833 31515 14867
rect 31549 14833 31587 14867
rect 31621 14833 31659 14867
rect 31693 14833 31731 14867
rect 31765 14833 31803 14867
rect 31837 14833 31875 14867
rect 31909 14833 31947 14867
rect 31981 14833 32019 14867
rect 32053 14833 32091 14867
rect 32125 14833 32163 14867
rect 32197 14833 32235 14867
rect 32269 14833 32307 14867
rect 32341 14833 32379 14867
rect 32413 14833 32451 14867
rect 32485 14833 32523 14867
rect 32557 14833 32595 14867
rect 32629 14833 32667 14867
rect 32701 14833 32739 14867
rect 32773 14833 32811 14867
rect 32845 14833 32883 14867
rect 32917 14833 32955 14867
rect 32989 14833 33027 14867
rect 33061 14833 33099 14867
rect 33133 14833 33171 14867
rect 33205 14833 33243 14867
rect 33277 14833 33315 14867
rect 33349 14833 33387 14867
rect 33421 14833 33459 14867
rect 33493 14833 33531 14867
rect 33565 14833 33603 14867
rect 33637 14833 33675 14867
rect 33709 14833 33747 14867
rect 33781 14833 33819 14867
rect 33853 14833 33891 14867
rect 33925 14833 33963 14867
rect 33997 14833 34035 14867
rect 34069 14833 34107 14867
rect 34141 14833 34179 14867
rect 34213 14833 34251 14867
rect 34285 14833 34323 14867
rect 34357 14833 34395 14867
rect 34429 14833 34467 14867
rect 34501 14833 34539 14867
rect 34573 14833 34611 14867
rect 34645 14833 34683 14867
rect 34717 14833 34755 14867
rect 34789 14833 34827 14867
rect 34861 14833 34899 14867
rect 34933 14833 34971 14867
rect 35005 14833 35043 14867
rect 35077 14833 35115 14867
rect 35149 14833 35187 14867
rect 35221 14833 35400 14867
rect -17500 14800 35400 14833
rect -17500 14797 -17400 14800
rect -17500 14763 -17467 14797
rect -17433 14763 -17400 14797
rect -17500 14725 -17400 14763
rect -17500 14691 -17467 14725
rect -17433 14691 -17400 14725
rect -17500 14653 -17400 14691
rect -17500 14619 -17467 14653
rect -17433 14619 -17400 14653
rect -17500 14581 -17400 14619
rect -17500 14547 -17467 14581
rect -17433 14547 -17400 14581
rect -17500 14509 -17400 14547
rect -17500 14475 -17467 14509
rect -17433 14475 -17400 14509
rect -17500 14437 -17400 14475
rect -17500 14403 -17467 14437
rect -17433 14403 -17400 14437
rect -17500 14365 -17400 14403
rect -17500 14331 -17467 14365
rect -17433 14331 -17400 14365
rect -17500 14293 -17400 14331
rect -17500 14259 -17467 14293
rect -17433 14259 -17400 14293
rect -17500 14221 -17400 14259
rect -17500 14187 -17467 14221
rect -17433 14187 -17400 14221
rect -17500 14149 -17400 14187
rect -17500 14115 -17467 14149
rect -17433 14115 -17400 14149
rect -17500 14077 -17400 14115
rect -17500 14043 -17467 14077
rect -17433 14043 -17400 14077
rect -17500 14005 -17400 14043
rect -17500 13971 -17467 14005
rect -17433 13971 -17400 14005
rect -17500 13933 -17400 13971
rect -17500 13899 -17467 13933
rect -17433 13899 -17400 13933
rect -17500 13861 -17400 13899
rect -17500 13827 -17467 13861
rect -17433 13827 -17400 13861
rect -17500 13789 -17400 13827
rect -17500 13755 -17467 13789
rect -17433 13755 -17400 13789
rect -17500 13717 -17400 13755
rect -17500 13683 -17467 13717
rect -17433 13683 -17400 13717
rect -17500 13645 -17400 13683
rect -17500 13611 -17467 13645
rect -17433 13611 -17400 13645
rect -17500 13573 -17400 13611
rect -17500 13539 -17467 13573
rect -17433 13539 -17400 13573
rect -17500 13501 -17400 13539
rect -17500 13467 -17467 13501
rect -17433 13467 -17400 13501
rect -17500 13429 -17400 13467
rect -17500 13395 -17467 13429
rect -17433 13395 -17400 13429
rect -17500 13357 -17400 13395
rect -17500 13323 -17467 13357
rect -17433 13323 -17400 13357
rect -17500 13285 -17400 13323
rect -17500 13251 -17467 13285
rect -17433 13251 -17400 13285
rect -17500 13213 -17400 13251
rect -17500 13179 -17467 13213
rect -17433 13179 -17400 13213
rect -17500 13141 -17400 13179
rect -17500 13107 -17467 13141
rect -17433 13107 -17400 13141
rect -17500 13069 -17400 13107
rect -17500 13035 -17467 13069
rect -17433 13035 -17400 13069
rect -17500 13020 -17400 13035
rect 35300 14797 35400 14800
rect 35300 14763 35333 14797
rect 35367 14763 35400 14797
rect 35300 14725 35400 14763
rect 35300 14691 35333 14725
rect 35367 14691 35400 14725
rect 35300 14653 35400 14691
rect 35300 14619 35333 14653
rect 35367 14619 35400 14653
rect 35300 14581 35400 14619
rect 35300 14547 35333 14581
rect 35367 14547 35400 14581
rect 35300 14509 35400 14547
rect 35300 14475 35333 14509
rect 35367 14475 35400 14509
rect 35300 14437 35400 14475
rect 35300 14403 35333 14437
rect 35367 14403 35400 14437
rect 35300 14365 35400 14403
rect 35300 14331 35333 14365
rect 35367 14331 35400 14365
rect 35300 14293 35400 14331
rect 35300 14259 35333 14293
rect 35367 14259 35400 14293
rect 35300 14221 35400 14259
rect 35300 14187 35333 14221
rect 35367 14187 35400 14221
rect 35300 14149 35400 14187
rect 35300 14115 35333 14149
rect 35367 14115 35400 14149
rect 35300 14077 35400 14115
rect 35300 14043 35333 14077
rect 35367 14043 35400 14077
rect 35300 14005 35400 14043
rect 35300 13971 35333 14005
rect 35367 13971 35400 14005
rect 35300 13933 35400 13971
rect 35300 13899 35333 13933
rect 35367 13899 35400 13933
rect 35300 13861 35400 13899
rect 35300 13827 35333 13861
rect 35367 13827 35400 13861
rect 35300 13789 35400 13827
rect 35300 13755 35333 13789
rect 35367 13755 35400 13789
rect 35300 13717 35400 13755
rect 35300 13683 35333 13717
rect 35367 13683 35400 13717
rect 35300 13645 35400 13683
rect 35300 13611 35333 13645
rect 35367 13611 35400 13645
rect 35300 13573 35400 13611
rect 35300 13539 35333 13573
rect 35367 13539 35400 13573
rect 35300 13501 35400 13539
rect 35300 13467 35333 13501
rect 35367 13467 35400 13501
rect 35300 13429 35400 13467
rect 35300 13395 35333 13429
rect 35367 13395 35400 13429
rect 35300 13357 35400 13395
rect 35300 13323 35333 13357
rect 35367 13323 35400 13357
rect 35300 13285 35400 13323
rect 35300 13251 35333 13285
rect 35367 13251 35400 13285
rect 35300 13213 35400 13251
rect 35300 13179 35333 13213
rect 35367 13179 35400 13213
rect 35300 13141 35400 13179
rect 35300 13107 35333 13141
rect 35367 13107 35400 13141
rect 35300 13069 35400 13107
rect 35300 13035 35333 13069
rect 35367 13035 35400 13069
rect 35300 13020 35400 13035
rect -17500 12997 35400 13020
rect -17500 12963 -17467 12997
rect -17433 12963 35333 12997
rect 35367 12963 35400 12997
rect -17500 12940 35400 12963
rect -17500 12925 -17400 12940
rect -17500 12891 -17467 12925
rect -17433 12891 -17400 12925
rect -17500 12853 -17400 12891
rect -17500 12819 -17467 12853
rect -17433 12819 -17400 12853
rect -17500 12781 -17400 12819
rect -17500 12747 -17467 12781
rect -17433 12747 -17400 12781
rect -17500 12709 -17400 12747
rect -17500 12675 -17467 12709
rect -17433 12675 -17400 12709
rect -17500 12637 -17400 12675
rect -17500 12603 -17467 12637
rect -17433 12603 -17400 12637
rect -17500 12565 -17400 12603
rect -17500 12531 -17467 12565
rect -17433 12531 -17400 12565
rect -17500 12493 -17400 12531
rect -17500 12459 -17467 12493
rect -17433 12459 -17400 12493
rect -17500 12421 -17400 12459
rect -17500 12387 -17467 12421
rect -17433 12387 -17400 12421
rect -17500 12349 -17400 12387
rect -17500 12315 -17467 12349
rect -17433 12315 -17400 12349
rect -17500 12277 -17400 12315
rect -17500 12243 -17467 12277
rect -17433 12243 -17400 12277
rect -17500 12205 -17400 12243
rect -17500 12171 -17467 12205
rect -17433 12171 -17400 12205
rect -17500 12133 -17400 12171
rect -17500 12099 -17467 12133
rect -17433 12099 -17400 12133
rect -17500 12061 -17400 12099
rect -17500 12027 -17467 12061
rect -17433 12027 -17400 12061
rect -17500 11989 -17400 12027
rect -17500 11955 -17467 11989
rect -17433 11955 -17400 11989
rect -17500 11917 -17400 11955
rect -17500 11883 -17467 11917
rect -17433 11883 -17400 11917
rect -17500 11845 -17400 11883
rect -17500 11811 -17467 11845
rect -17433 11811 -17400 11845
rect -17500 11773 -17400 11811
rect -17500 11739 -17467 11773
rect -17433 11739 -17400 11773
rect -17500 11701 -17400 11739
rect -17500 11667 -17467 11701
rect -17433 11667 -17400 11701
rect -17500 11629 -17400 11667
rect -17500 11595 -17467 11629
rect -17433 11595 -17400 11629
rect -17500 11557 -17400 11595
rect -17500 11523 -17467 11557
rect -17433 11523 -17400 11557
rect -17500 11485 -17400 11523
rect -17500 11451 -17467 11485
rect -17433 11451 -17400 11485
rect -17500 11413 -17400 11451
rect -17500 11379 -17467 11413
rect -17433 11379 -17400 11413
rect -17500 11341 -17400 11379
rect -17500 11307 -17467 11341
rect -17433 11307 -17400 11341
rect -17500 11269 -17400 11307
rect -17500 11235 -17467 11269
rect -17433 11235 -17400 11269
rect -17500 11197 -17400 11235
rect -17500 11163 -17467 11197
rect -17433 11163 -17400 11197
rect -17500 11125 -17400 11163
rect -17500 11091 -17467 11125
rect -17433 11091 -17400 11125
rect -17500 11053 -17400 11091
rect -17500 11019 -17467 11053
rect -17433 11019 -17400 11053
rect -17500 10981 -17400 11019
rect -17500 10947 -17467 10981
rect -17433 10947 -17400 10981
rect -17500 10909 -17400 10947
rect -17500 10875 -17467 10909
rect -17433 10875 -17400 10909
rect -17500 10837 -17400 10875
rect -17500 10803 -17467 10837
rect -17433 10803 -17400 10837
rect -17500 10765 -17400 10803
rect -17500 10731 -17467 10765
rect -17433 10731 -17400 10765
rect -17500 10693 -17400 10731
rect -17500 10659 -17467 10693
rect -17433 10659 -17400 10693
rect -17500 10621 -17400 10659
rect -17500 10587 -17467 10621
rect -17433 10587 -17400 10621
rect -17500 10549 -17400 10587
rect -17500 10515 -17467 10549
rect -17433 10515 -17400 10549
rect -17500 10477 -17400 10515
rect -17500 10443 -17467 10477
rect -17433 10443 -17400 10477
rect -17500 10405 -17400 10443
rect -17500 10371 -17467 10405
rect -17433 10371 -17400 10405
rect -17500 10333 -17400 10371
rect -17500 10299 -17467 10333
rect -17433 10299 -17400 10333
rect -17500 10261 -17400 10299
rect -17500 10227 -17467 10261
rect -17433 10227 -17400 10261
rect -17500 10189 -17400 10227
rect -17500 10155 -17467 10189
rect -17433 10155 -17400 10189
rect -17500 10117 -17400 10155
rect -17500 10083 -17467 10117
rect -17433 10083 -17400 10117
rect -17500 10045 -17400 10083
rect -17500 10011 -17467 10045
rect -17433 10011 -17400 10045
rect -17500 9973 -17400 10011
rect -17500 9939 -17467 9973
rect -17433 9939 -17400 9973
rect -17500 9901 -17400 9939
rect -17500 9867 -17467 9901
rect -17433 9867 -17400 9901
rect -17500 9829 -17400 9867
rect -17500 9795 -17467 9829
rect -17433 9795 -17400 9829
rect -17500 9757 -17400 9795
rect -17500 9723 -17467 9757
rect -17433 9723 -17400 9757
rect -17500 9685 -17400 9723
rect -17500 9651 -17467 9685
rect -17433 9651 -17400 9685
rect -17500 9613 -17400 9651
rect -17500 9579 -17467 9613
rect -17433 9579 -17400 9613
rect -17500 9541 -17400 9579
rect -17500 9507 -17467 9541
rect -17433 9507 -17400 9541
rect -17500 9500 -17400 9507
rect 35300 12925 35400 12940
rect 35300 12891 35333 12925
rect 35367 12891 35400 12925
rect 35300 12853 35400 12891
rect 35300 12819 35333 12853
rect 35367 12819 35400 12853
rect 35300 12781 35400 12819
rect 35300 12747 35333 12781
rect 35367 12747 35400 12781
rect 35300 12709 35400 12747
rect 35300 12675 35333 12709
rect 35367 12675 35400 12709
rect 35300 12637 35400 12675
rect 35300 12603 35333 12637
rect 35367 12603 35400 12637
rect 35300 12565 35400 12603
rect 35300 12531 35333 12565
rect 35367 12531 35400 12565
rect 35300 12493 35400 12531
rect 35300 12459 35333 12493
rect 35367 12459 35400 12493
rect 35300 12421 35400 12459
rect 35300 12387 35333 12421
rect 35367 12387 35400 12421
rect 35300 12349 35400 12387
rect 35300 12315 35333 12349
rect 35367 12315 35400 12349
rect 35300 12277 35400 12315
rect 35300 12243 35333 12277
rect 35367 12243 35400 12277
rect 35300 12205 35400 12243
rect 35300 12171 35333 12205
rect 35367 12171 35400 12205
rect 35300 12133 35400 12171
rect 35300 12099 35333 12133
rect 35367 12099 35400 12133
rect 35300 12061 35400 12099
rect 35300 12027 35333 12061
rect 35367 12027 35400 12061
rect 35300 11989 35400 12027
rect 35300 11955 35333 11989
rect 35367 11955 35400 11989
rect 35300 11917 35400 11955
rect 35300 11883 35333 11917
rect 35367 11883 35400 11917
rect 35300 11845 35400 11883
rect 35300 11811 35333 11845
rect 35367 11811 35400 11845
rect 35300 11773 35400 11811
rect 35300 11739 35333 11773
rect 35367 11739 35400 11773
rect 35300 11701 35400 11739
rect 35300 11667 35333 11701
rect 35367 11667 35400 11701
rect 35300 11629 35400 11667
rect 35300 11595 35333 11629
rect 35367 11595 35400 11629
rect 35300 11557 35400 11595
rect 35300 11523 35333 11557
rect 35367 11523 35400 11557
rect 35300 11485 35400 11523
rect 35300 11451 35333 11485
rect 35367 11451 35400 11485
rect 35300 11413 35400 11451
rect 35300 11379 35333 11413
rect 35367 11379 35400 11413
rect 35300 11341 35400 11379
rect 35300 11307 35333 11341
rect 35367 11307 35400 11341
rect 35300 11269 35400 11307
rect 35300 11235 35333 11269
rect 35367 11235 35400 11269
rect 35300 11197 35400 11235
rect 35300 11163 35333 11197
rect 35367 11163 35400 11197
rect 35300 11125 35400 11163
rect 35300 11091 35333 11125
rect 35367 11091 35400 11125
rect 35300 11053 35400 11091
rect 35300 11019 35333 11053
rect 35367 11019 35400 11053
rect 35300 10981 35400 11019
rect 35300 10947 35333 10981
rect 35367 10947 35400 10981
rect 35300 10909 35400 10947
rect 35300 10875 35333 10909
rect 35367 10875 35400 10909
rect 35300 10837 35400 10875
rect 35300 10803 35333 10837
rect 35367 10803 35400 10837
rect 35300 10765 35400 10803
rect 35300 10731 35333 10765
rect 35367 10731 35400 10765
rect 35300 10693 35400 10731
rect 35300 10659 35333 10693
rect 35367 10659 35400 10693
rect 35300 10621 35400 10659
rect 35300 10587 35333 10621
rect 35367 10587 35400 10621
rect 35300 10549 35400 10587
rect 35300 10515 35333 10549
rect 35367 10515 35400 10549
rect 35300 10477 35400 10515
rect 35300 10443 35333 10477
rect 35367 10443 35400 10477
rect 35300 10405 35400 10443
rect 35300 10371 35333 10405
rect 35367 10371 35400 10405
rect 35300 10333 35400 10371
rect 35300 10299 35333 10333
rect 35367 10299 35400 10333
rect 35300 10261 35400 10299
rect 35300 10227 35333 10261
rect 35367 10227 35400 10261
rect 35300 10189 35400 10227
rect 35300 10155 35333 10189
rect 35367 10155 35400 10189
rect 35300 10117 35400 10155
rect 35300 10083 35333 10117
rect 35367 10083 35400 10117
rect 35300 10045 35400 10083
rect 35300 10011 35333 10045
rect 35367 10011 35400 10045
rect 35300 9973 35400 10011
rect 35300 9939 35333 9973
rect 35367 9939 35400 9973
rect 35300 9901 35400 9939
rect 35300 9867 35333 9901
rect 35367 9867 35400 9901
rect 35300 9829 35400 9867
rect 35300 9795 35333 9829
rect 35367 9795 35400 9829
rect 35300 9757 35400 9795
rect 35300 9723 35333 9757
rect 35367 9723 35400 9757
rect 35300 9685 35400 9723
rect 35300 9651 35333 9685
rect 35367 9651 35400 9685
rect 35300 9613 35400 9651
rect 35300 9579 35333 9613
rect 35367 9579 35400 9613
rect 35300 9541 35400 9579
rect 35300 9507 35333 9541
rect 35367 9507 35400 9541
rect 35300 9500 35400 9507
rect -17500 9469 35400 9500
rect -17500 9435 -17467 9469
rect -17433 9435 35333 9469
rect 35367 9435 35400 9469
rect -17500 9420 35400 9435
rect -17500 9397 -17400 9420
rect -17500 9363 -17467 9397
rect -17433 9363 -17400 9397
rect -17500 9325 -17400 9363
rect -17500 9291 -17467 9325
rect -17433 9291 -17400 9325
rect -17500 9253 -17400 9291
rect -17500 9219 -17467 9253
rect -17433 9219 -17400 9253
rect -17500 9181 -17400 9219
rect -17500 9147 -17467 9181
rect -17433 9147 -17400 9181
rect -17500 9109 -17400 9147
rect -17500 9075 -17467 9109
rect -17433 9075 -17400 9109
rect -17500 9037 -17400 9075
rect -17500 9003 -17467 9037
rect -17433 9003 -17400 9037
rect -17500 8965 -17400 9003
rect -17500 8931 -17467 8965
rect -17433 8931 -17400 8965
rect -17500 8893 -17400 8931
rect -17500 8859 -17467 8893
rect -17433 8859 -17400 8893
rect -17500 8821 -17400 8859
rect -17500 8787 -17467 8821
rect -17433 8787 -17400 8821
rect -17500 8749 -17400 8787
rect -17500 8715 -17467 8749
rect -17433 8715 -17400 8749
rect -17500 8677 -17400 8715
rect -17500 8643 -17467 8677
rect -17433 8643 -17400 8677
rect -17500 8605 -17400 8643
rect -17500 8571 -17467 8605
rect -17433 8571 -17400 8605
rect -17500 8533 -17400 8571
rect -17500 8499 -17467 8533
rect -17433 8499 -17400 8533
rect -17500 8461 -17400 8499
rect -17500 8427 -17467 8461
rect -17433 8427 -17400 8461
rect -17500 8389 -17400 8427
rect -17500 8355 -17467 8389
rect -17433 8355 -17400 8389
rect -17500 8317 -17400 8355
rect -17500 8283 -17467 8317
rect -17433 8283 -17400 8317
rect -17500 8245 -17400 8283
rect -17500 8211 -17467 8245
rect -17433 8211 -17400 8245
rect -17500 8173 -17400 8211
rect -17500 8139 -17467 8173
rect -17433 8139 -17400 8173
rect -17500 8101 -17400 8139
rect -17500 8067 -17467 8101
rect -17433 8067 -17400 8101
rect -17500 8029 -17400 8067
rect -17500 7995 -17467 8029
rect -17433 7995 -17400 8029
rect -17500 7957 -17400 7995
rect -17500 7923 -17467 7957
rect -17433 7923 -17400 7957
rect -17500 7885 -17400 7923
rect -17500 7851 -17467 7885
rect -17433 7851 -17400 7885
rect -17500 7813 -17400 7851
rect -17500 7779 -17467 7813
rect -17433 7779 -17400 7813
rect -17500 7741 -17400 7779
rect -17500 7707 -17467 7741
rect -17433 7707 -17400 7741
rect -17500 7669 -17400 7707
rect -17500 7635 -17467 7669
rect -17433 7635 -17400 7669
rect -17500 7597 -17400 7635
rect -17500 7563 -17467 7597
rect -17433 7563 -17400 7597
rect -17500 7525 -17400 7563
rect -17500 7491 -17467 7525
rect -17433 7491 -17400 7525
rect -17500 7453 -17400 7491
rect -17500 7419 -17467 7453
rect -17433 7419 -17400 7453
rect -17500 7381 -17400 7419
rect -17500 7347 -17467 7381
rect -17433 7347 -17400 7381
rect -17500 7309 -17400 7347
rect -17500 7275 -17467 7309
rect -17433 7275 -17400 7309
rect -17500 7237 -17400 7275
rect -17500 7203 -17467 7237
rect -17433 7203 -17400 7237
rect -17500 7165 -17400 7203
rect -17500 7131 -17467 7165
rect -17433 7131 -17400 7165
rect -17500 7093 -17400 7131
rect -17500 7059 -17467 7093
rect -17433 7059 -17400 7093
rect -17500 7021 -17400 7059
rect -17500 6987 -17467 7021
rect -17433 6987 -17400 7021
rect -17500 6949 -17400 6987
rect -17500 6915 -17467 6949
rect -17433 6915 -17400 6949
rect -17500 6877 -17400 6915
rect -17500 6843 -17467 6877
rect -17433 6843 -17400 6877
rect -17500 6805 -17400 6843
rect -17500 6771 -17467 6805
rect -17433 6771 -17400 6805
rect -17500 6733 -17400 6771
rect -17500 6699 -17467 6733
rect -17433 6699 -17400 6733
rect -17500 6661 -17400 6699
rect -17500 6627 -17467 6661
rect -17433 6627 -17400 6661
rect -17500 6589 -17400 6627
rect -17500 6555 -17467 6589
rect -17433 6555 -17400 6589
rect -17500 6517 -17400 6555
rect -17500 6483 -17467 6517
rect -17433 6483 -17400 6517
rect -17500 6445 -17400 6483
rect -17500 6411 -17467 6445
rect -17433 6411 -17400 6445
rect -17500 6373 -17400 6411
rect -17500 6339 -17467 6373
rect -17433 6339 -17400 6373
rect -17500 6301 -17400 6339
rect -17500 6267 -17467 6301
rect -17433 6267 -17400 6301
rect -17500 6229 -17400 6267
rect -17500 6195 -17467 6229
rect -17433 6195 -17400 6229
rect -17500 6157 -17400 6195
rect -17500 6123 -17467 6157
rect -17433 6123 -17400 6157
rect -17500 6085 -17400 6123
rect -17500 6051 -17467 6085
rect -17433 6051 -17400 6085
rect -17500 6013 -17400 6051
rect -17500 5979 -17467 6013
rect -17433 5979 -17400 6013
rect -17500 5941 -17400 5979
rect -17500 5907 -17467 5941
rect -17433 5907 -17400 5941
rect -17500 5869 -17400 5907
rect -17500 5835 -17467 5869
rect -17433 5835 -17400 5869
rect -17500 5797 -17400 5835
rect -17500 5763 -17467 5797
rect -17433 5763 -17400 5797
rect -17500 5725 -17400 5763
rect 35300 9397 35400 9420
rect 35300 9363 35333 9397
rect 35367 9363 35400 9397
rect 35300 9325 35400 9363
rect 35300 9291 35333 9325
rect 35367 9291 35400 9325
rect 35300 9253 35400 9291
rect 35300 9219 35333 9253
rect 35367 9219 35400 9253
rect 35300 9181 35400 9219
rect 35300 9147 35333 9181
rect 35367 9147 35400 9181
rect 35300 9109 35400 9147
rect 35300 9075 35333 9109
rect 35367 9075 35400 9109
rect 35300 9037 35400 9075
rect 35300 9003 35333 9037
rect 35367 9003 35400 9037
rect 35300 8965 35400 9003
rect 35300 8931 35333 8965
rect 35367 8931 35400 8965
rect 35300 8893 35400 8931
rect 35300 8859 35333 8893
rect 35367 8859 35400 8893
rect 35300 8821 35400 8859
rect 35300 8787 35333 8821
rect 35367 8787 35400 8821
rect 35300 8749 35400 8787
rect 35300 8715 35333 8749
rect 35367 8715 35400 8749
rect 35300 8677 35400 8715
rect 35300 8643 35333 8677
rect 35367 8643 35400 8677
rect 35300 8605 35400 8643
rect 35300 8571 35333 8605
rect 35367 8571 35400 8605
rect 35300 8533 35400 8571
rect 35300 8499 35333 8533
rect 35367 8499 35400 8533
rect 35300 8461 35400 8499
rect 35300 8427 35333 8461
rect 35367 8427 35400 8461
rect 35300 8389 35400 8427
rect 35300 8355 35333 8389
rect 35367 8355 35400 8389
rect 35300 8317 35400 8355
rect 35300 8283 35333 8317
rect 35367 8283 35400 8317
rect 35300 8245 35400 8283
rect 35300 8211 35333 8245
rect 35367 8211 35400 8245
rect 35300 8173 35400 8211
rect 35300 8139 35333 8173
rect 35367 8139 35400 8173
rect 35300 8101 35400 8139
rect 35300 8067 35333 8101
rect 35367 8067 35400 8101
rect 35300 8029 35400 8067
rect 35300 7995 35333 8029
rect 35367 7995 35400 8029
rect 35300 7957 35400 7995
rect 35300 7923 35333 7957
rect 35367 7923 35400 7957
rect 35300 7885 35400 7923
rect 35300 7851 35333 7885
rect 35367 7851 35400 7885
rect 35300 7813 35400 7851
rect 35300 7779 35333 7813
rect 35367 7779 35400 7813
rect 35300 7741 35400 7779
rect 35300 7707 35333 7741
rect 35367 7707 35400 7741
rect 35300 7669 35400 7707
rect 35300 7635 35333 7669
rect 35367 7635 35400 7669
rect 35300 7597 35400 7635
rect 35300 7563 35333 7597
rect 35367 7563 35400 7597
rect 35300 7525 35400 7563
rect 35300 7491 35333 7525
rect 35367 7491 35400 7525
rect 35300 7453 35400 7491
rect 35300 7419 35333 7453
rect 35367 7419 35400 7453
rect 35300 7381 35400 7419
rect 35300 7347 35333 7381
rect 35367 7347 35400 7381
rect 35300 7309 35400 7347
rect 35300 7275 35333 7309
rect 35367 7275 35400 7309
rect 35300 7237 35400 7275
rect 35300 7203 35333 7237
rect 35367 7203 35400 7237
rect 35300 7165 35400 7203
rect 35300 7131 35333 7165
rect 35367 7131 35400 7165
rect 35300 7093 35400 7131
rect 35300 7059 35333 7093
rect 35367 7059 35400 7093
rect 35300 7021 35400 7059
rect 35300 6987 35333 7021
rect 35367 6987 35400 7021
rect 35300 6949 35400 6987
rect 35300 6915 35333 6949
rect 35367 6915 35400 6949
rect 35300 6877 35400 6915
rect 35300 6843 35333 6877
rect 35367 6843 35400 6877
rect 35300 6805 35400 6843
rect 35300 6771 35333 6805
rect 35367 6771 35400 6805
rect 35300 6733 35400 6771
rect 35300 6699 35333 6733
rect 35367 6699 35400 6733
rect 35300 6661 35400 6699
rect 35300 6627 35333 6661
rect 35367 6627 35400 6661
rect 35300 6589 35400 6627
rect 35300 6555 35333 6589
rect 35367 6555 35400 6589
rect 35300 6517 35400 6555
rect 35300 6483 35333 6517
rect 35367 6483 35400 6517
rect 35300 6445 35400 6483
rect 35300 6411 35333 6445
rect 35367 6411 35400 6445
rect 35300 6373 35400 6411
rect 35300 6339 35333 6373
rect 35367 6339 35400 6373
rect 35300 6301 35400 6339
rect 35300 6267 35333 6301
rect 35367 6267 35400 6301
rect 35300 6229 35400 6267
rect 35300 6195 35333 6229
rect 35367 6195 35400 6229
rect 35300 6157 35400 6195
rect 35300 6123 35333 6157
rect 35367 6123 35400 6157
rect 35300 6085 35400 6123
rect 35300 6051 35333 6085
rect 35367 6051 35400 6085
rect 35300 6013 35400 6051
rect 35300 5979 35333 6013
rect 35367 5979 35400 6013
rect 35300 5941 35400 5979
rect 35300 5907 35333 5941
rect 35367 5907 35400 5941
rect 35300 5869 35400 5907
rect 35300 5835 35333 5869
rect 35367 5835 35400 5869
rect 35300 5797 35400 5835
rect 35300 5763 35333 5797
rect 35367 5763 35400 5797
rect -17500 5691 -17467 5725
rect -17433 5691 -17400 5725
rect -17500 5653 -17400 5691
rect -17500 5619 -17467 5653
rect -17433 5620 -17400 5653
rect -17433 5619 200 5620
rect -17500 5581 200 5619
rect -17500 5547 -17467 5581
rect -17433 5547 200 5581
rect -17500 5540 200 5547
rect -17500 5509 -17400 5540
rect -17500 5475 -17467 5509
rect -17433 5475 -17400 5509
rect -17500 5437 -17400 5475
rect -17500 5403 -17467 5437
rect -17433 5403 -17400 5437
rect 300 5420 420 5740
rect 2060 5640 2180 5740
rect 35300 5725 35400 5763
rect 35300 5691 35333 5725
rect 35367 5691 35400 5725
rect 35300 5653 35400 5691
rect 2060 5520 2600 5640
rect 4280 5520 4800 5640
rect 6480 5520 7000 5640
rect 8680 5520 9200 5640
rect 10880 5520 11400 5640
rect 13080 5520 13600 5640
rect 15280 5520 15800 5640
rect 35300 5620 35333 5653
rect 17780 5619 35333 5620
rect 35367 5619 35400 5653
rect 17780 5581 35400 5619
rect 17780 5547 35333 5581
rect 35367 5547 35400 5581
rect 17780 5540 35400 5547
rect 2060 5420 2180 5520
rect 35300 5509 35400 5540
rect 35300 5475 35333 5509
rect 35367 5475 35400 5509
rect 35300 5437 35400 5475
rect -17500 5365 -17400 5403
rect -17500 5331 -17467 5365
rect -17433 5331 -17400 5365
rect -17500 5293 -17400 5331
rect -17500 5259 -17467 5293
rect -17433 5259 -17400 5293
rect -17500 5221 -17400 5259
rect -17500 5187 -17467 5221
rect -17433 5187 -17400 5221
rect -17500 5149 -17400 5187
rect -17500 5115 -17467 5149
rect -17433 5115 -17400 5149
rect -17500 5077 -17400 5115
rect -17500 5043 -17467 5077
rect -17433 5043 -17400 5077
rect -17500 5005 -17400 5043
rect -17500 4971 -17467 5005
rect -17433 4971 -17400 5005
rect -17500 4933 -17400 4971
rect -17500 4899 -17467 4933
rect -17433 4899 -17400 4933
rect -17500 4861 -17400 4899
rect -17500 4827 -17467 4861
rect -17433 4827 -17400 4861
rect -17500 4789 -17400 4827
rect -17500 4755 -17467 4789
rect -17433 4755 -17400 4789
rect -17500 4717 -17400 4755
rect -17500 4683 -17467 4717
rect -17433 4683 -17400 4717
rect -17500 4645 -17400 4683
rect -17500 4611 -17467 4645
rect -17433 4611 -17400 4645
rect -17500 4573 -17400 4611
rect -17500 4539 -17467 4573
rect -17433 4539 -17400 4573
rect -17500 4501 -17400 4539
rect -17500 4467 -17467 4501
rect -17433 4467 -17400 4501
rect -17500 4429 -17400 4467
rect -17500 4395 -17467 4429
rect -17433 4395 -17400 4429
rect -17500 4357 -17400 4395
rect -17500 4323 -17467 4357
rect -17433 4323 -17400 4357
rect -17500 4285 -17400 4323
rect -17500 4251 -17467 4285
rect -17433 4251 -17400 4285
rect -17500 4213 -17400 4251
rect -17500 4179 -17467 4213
rect -17433 4179 -17400 4213
rect -17500 4141 -17400 4179
rect -17500 4107 -17467 4141
rect -17433 4107 -17400 4141
rect -17500 4069 -17400 4107
rect -17500 4035 -17467 4069
rect -17433 4035 -17400 4069
rect -17500 3997 -17400 4035
rect -17500 3963 -17467 3997
rect -17433 3963 -17400 3997
rect -17500 3925 -17400 3963
rect -17500 3891 -17467 3925
rect -17433 3891 -17400 3925
rect -17500 3853 -17400 3891
rect -17500 3819 -17467 3853
rect -17433 3819 -17400 3853
rect -17500 3781 -17400 3819
rect -17500 3747 -17467 3781
rect -17433 3747 -17400 3781
rect -17500 3709 -17400 3747
rect -17500 3675 -17467 3709
rect -17433 3675 -17400 3709
rect -17500 3637 -17400 3675
rect -17500 3603 -17467 3637
rect -17433 3603 -17400 3637
rect -17500 3565 -17400 3603
rect -17500 3531 -17467 3565
rect -17433 3531 -17400 3565
rect -17500 3493 -17400 3531
rect -17500 3459 -17467 3493
rect -17433 3459 -17400 3493
rect -17500 3421 -17400 3459
rect -17500 3387 -17467 3421
rect -17433 3387 -17400 3421
rect -17500 3349 -17400 3387
rect -17500 3315 -17467 3349
rect -17433 3315 -17400 3349
rect -17500 3277 -17400 3315
rect -17500 3243 -17467 3277
rect -17433 3243 -17400 3277
rect -17500 3205 -17400 3243
rect -17500 3171 -17467 3205
rect -17433 3171 -17400 3205
rect -17500 3133 -17400 3171
rect -17500 3099 -17467 3133
rect -17433 3099 -17400 3133
rect -17500 3061 -17400 3099
rect -17500 3027 -17467 3061
rect -17433 3027 -17400 3061
rect -17500 2989 -17400 3027
rect -17500 2955 -17467 2989
rect -17433 2955 -17400 2989
rect -17500 2917 -17400 2955
rect -17500 2883 -17467 2917
rect -17433 2883 -17400 2917
rect -17500 2845 -17400 2883
rect -17500 2811 -17467 2845
rect -17433 2811 -17400 2845
rect -17500 2773 -17400 2811
rect -17500 2739 -17467 2773
rect -17433 2739 -17400 2773
rect -17500 2701 -17400 2739
rect -17500 2667 -17467 2701
rect -17433 2667 -17400 2701
rect -17500 2629 -17400 2667
rect -17500 2595 -17467 2629
rect -17433 2595 -17400 2629
rect -17500 2557 -17400 2595
rect -17500 2523 -17467 2557
rect -17433 2523 -17400 2557
rect -17500 2485 -17400 2523
rect -17500 2451 -17467 2485
rect -17433 2451 -17400 2485
rect -17500 2413 -17400 2451
rect -17500 2379 -17467 2413
rect -17433 2379 -17400 2413
rect -17500 2341 -17400 2379
rect -17500 2307 -17467 2341
rect -17433 2307 -17400 2341
rect -17500 2269 -17400 2307
rect -17500 2235 -17467 2269
rect -17433 2235 -17400 2269
rect -17500 2197 -17400 2235
rect 35300 5403 35333 5437
rect 35367 5403 35400 5437
rect 35300 5365 35400 5403
rect 35300 5331 35333 5365
rect 35367 5331 35400 5365
rect 35300 5293 35400 5331
rect 35300 5259 35333 5293
rect 35367 5259 35400 5293
rect 35300 5221 35400 5259
rect 35300 5187 35333 5221
rect 35367 5187 35400 5221
rect 35300 5149 35400 5187
rect 35300 5115 35333 5149
rect 35367 5115 35400 5149
rect 35300 5077 35400 5115
rect 35300 5043 35333 5077
rect 35367 5043 35400 5077
rect 35300 5005 35400 5043
rect 35300 4971 35333 5005
rect 35367 4971 35400 5005
rect 35300 4933 35400 4971
rect 35300 4899 35333 4933
rect 35367 4899 35400 4933
rect 35300 4861 35400 4899
rect 35300 4827 35333 4861
rect 35367 4827 35400 4861
rect 35300 4789 35400 4827
rect 35300 4755 35333 4789
rect 35367 4755 35400 4789
rect 35300 4717 35400 4755
rect 35300 4683 35333 4717
rect 35367 4683 35400 4717
rect 35300 4645 35400 4683
rect 35300 4611 35333 4645
rect 35367 4611 35400 4645
rect 35300 4573 35400 4611
rect 35300 4539 35333 4573
rect 35367 4539 35400 4573
rect 35300 4501 35400 4539
rect 35300 4467 35333 4501
rect 35367 4467 35400 4501
rect 35300 4429 35400 4467
rect 35300 4395 35333 4429
rect 35367 4395 35400 4429
rect 35300 4357 35400 4395
rect 35300 4323 35333 4357
rect 35367 4323 35400 4357
rect 35300 4285 35400 4323
rect 35300 4251 35333 4285
rect 35367 4251 35400 4285
rect 35300 4213 35400 4251
rect 35300 4179 35333 4213
rect 35367 4179 35400 4213
rect 35300 4141 35400 4179
rect 35300 4107 35333 4141
rect 35367 4107 35400 4141
rect 35300 4069 35400 4107
rect 35300 4035 35333 4069
rect 35367 4035 35400 4069
rect 35300 3997 35400 4035
rect 35300 3963 35333 3997
rect 35367 3963 35400 3997
rect 35300 3925 35400 3963
rect 35300 3891 35333 3925
rect 35367 3891 35400 3925
rect 35300 3853 35400 3891
rect 35300 3819 35333 3853
rect 35367 3819 35400 3853
rect 35300 3781 35400 3819
rect 35300 3747 35333 3781
rect 35367 3747 35400 3781
rect 35300 3709 35400 3747
rect 35300 3675 35333 3709
rect 35367 3675 35400 3709
rect 35300 3637 35400 3675
rect 35300 3603 35333 3637
rect 35367 3603 35400 3637
rect 35300 3565 35400 3603
rect 35300 3531 35333 3565
rect 35367 3531 35400 3565
rect 35300 3493 35400 3531
rect 35300 3459 35333 3493
rect 35367 3459 35400 3493
rect 35300 3421 35400 3459
rect 35300 3387 35333 3421
rect 35367 3387 35400 3421
rect 35300 3349 35400 3387
rect 35300 3315 35333 3349
rect 35367 3315 35400 3349
rect 35300 3277 35400 3315
rect 35300 3243 35333 3277
rect 35367 3243 35400 3277
rect 35300 3205 35400 3243
rect 35300 3171 35333 3205
rect 35367 3171 35400 3205
rect 35300 3133 35400 3171
rect 35300 3099 35333 3133
rect 35367 3099 35400 3133
rect 35300 3061 35400 3099
rect 35300 3027 35333 3061
rect 35367 3027 35400 3061
rect 35300 2989 35400 3027
rect 35300 2955 35333 2989
rect 35367 2955 35400 2989
rect 35300 2917 35400 2955
rect 35300 2883 35333 2917
rect 35367 2883 35400 2917
rect 35300 2845 35400 2883
rect 35300 2811 35333 2845
rect 35367 2811 35400 2845
rect 35300 2773 35400 2811
rect 35300 2739 35333 2773
rect 35367 2739 35400 2773
rect 35300 2701 35400 2739
rect 35300 2667 35333 2701
rect 35367 2667 35400 2701
rect 35300 2629 35400 2667
rect 35300 2595 35333 2629
rect 35367 2595 35400 2629
rect 35300 2557 35400 2595
rect 35300 2523 35333 2557
rect 35367 2523 35400 2557
rect 35300 2485 35400 2523
rect 35300 2451 35333 2485
rect 35367 2451 35400 2485
rect 35300 2413 35400 2451
rect 35300 2379 35333 2413
rect 35367 2379 35400 2413
rect 35300 2341 35400 2379
rect 35300 2307 35333 2341
rect 35367 2307 35400 2341
rect 35300 2269 35400 2307
rect 35300 2235 35333 2269
rect 35367 2235 35400 2269
rect -17500 2163 -17467 2197
rect -17433 2163 -17400 2197
rect -17500 2125 -17400 2163
rect -17500 2091 -17467 2125
rect -17433 2100 -17400 2125
rect -17433 2091 200 2100
rect -17500 2053 200 2091
rect -17500 2019 -17467 2053
rect -17433 2020 200 2053
rect -17433 2019 -17400 2020
rect -17500 1981 -17400 2019
rect -17500 1947 -17467 1981
rect -17433 1947 -17400 1981
rect -17500 1909 -17400 1947
rect 740 1920 840 2200
rect 1660 1940 1760 2220
rect 35300 2197 35400 2235
rect 35300 2163 35333 2197
rect 35367 2163 35400 2197
rect 35300 2125 35400 2163
rect 2080 2020 2620 2120
rect 4260 2020 4800 2120
rect 6460 2020 7000 2120
rect 8680 2020 9220 2120
rect 10880 2020 11420 2120
rect 13060 2020 13600 2120
rect 15280 2020 15820 2120
rect 35300 2100 35333 2125
rect 17780 2091 35333 2100
rect 35367 2091 35400 2125
rect 17780 2053 35400 2091
rect 17780 2020 35333 2053
rect 35300 2019 35333 2020
rect 35367 2019 35400 2053
rect 35300 1981 35400 2019
rect 35300 1947 35333 1981
rect 35367 1947 35400 1981
rect -17500 1875 -17467 1909
rect -17433 1875 -17400 1909
rect -17500 1837 -17400 1875
rect -17500 1803 -17467 1837
rect -17433 1803 -17400 1837
rect -17500 1765 -17400 1803
rect -17500 1731 -17467 1765
rect -17433 1731 -17400 1765
rect -17500 1693 -17400 1731
rect -17500 1659 -17467 1693
rect -17433 1659 -17400 1693
rect -17500 1621 -17400 1659
rect -17500 1587 -17467 1621
rect -17433 1587 -17400 1621
rect -17500 1549 -17400 1587
rect -17500 1515 -17467 1549
rect -17433 1515 -17400 1549
rect -17500 1477 -17400 1515
rect -17500 1443 -17467 1477
rect -17433 1443 -17400 1477
rect -17500 1405 -17400 1443
rect -17500 1371 -17467 1405
rect -17433 1371 -17400 1405
rect -17500 1333 -17400 1371
rect -17500 1299 -17467 1333
rect -17433 1299 -17400 1333
rect -17500 1261 -17400 1299
rect -17500 1227 -17467 1261
rect -17433 1227 -17400 1261
rect -17500 1189 -17400 1227
rect -17500 1155 -17467 1189
rect -17433 1155 -17400 1189
rect -17500 1117 -17400 1155
rect -17500 1083 -17467 1117
rect -17433 1083 -17400 1117
rect -17500 1045 -17400 1083
rect -17500 1011 -17467 1045
rect -17433 1011 -17400 1045
rect -17500 973 -17400 1011
rect -17500 939 -17467 973
rect -17433 939 -17400 973
rect -17500 901 -17400 939
rect -17500 867 -17467 901
rect -17433 867 -17400 901
rect -17500 829 -17400 867
rect -17500 795 -17467 829
rect -17433 795 -17400 829
rect -17500 757 -17400 795
rect -17500 723 -17467 757
rect -17433 723 -17400 757
rect -17500 685 -17400 723
rect -17500 651 -17467 685
rect -17433 651 -17400 685
rect -17500 613 -17400 651
rect -17500 579 -17467 613
rect -17433 579 -17400 613
rect -17500 541 -17400 579
rect -17500 507 -17467 541
rect -17433 507 -17400 541
rect -17500 469 -17400 507
rect -17500 435 -17467 469
rect -17433 435 -17400 469
rect -17500 397 -17400 435
rect -17500 363 -17467 397
rect -17433 363 -17400 397
rect -17500 325 -17400 363
rect -17500 291 -17467 325
rect -17433 291 -17400 325
rect -17500 253 -17400 291
rect -17500 219 -17467 253
rect -17433 219 -17400 253
rect -17500 181 -17400 219
rect -17500 147 -17467 181
rect -17433 147 -17400 181
rect -17500 109 -17400 147
rect -17500 75 -17467 109
rect -17433 75 -17400 109
rect -17500 37 -17400 75
rect -17500 3 -17467 37
rect -17433 3 -17400 37
rect -17500 -35 -17400 3
rect -17500 -69 -17467 -35
rect -17433 -69 -17400 -35
rect -17500 -107 -17400 -69
rect -17500 -141 -17467 -107
rect -17433 -141 -17400 -107
rect -17500 -179 -17400 -141
rect -17500 -213 -17467 -179
rect -17433 -213 -17400 -179
rect -17500 -251 -17400 -213
rect -17500 -285 -17467 -251
rect -17433 -285 -17400 -251
rect -17500 -323 -17400 -285
rect -17500 -357 -17467 -323
rect -17433 -357 -17400 -323
rect -17500 -395 -17400 -357
rect -17500 -429 -17467 -395
rect -17433 -429 -17400 -395
rect -17500 -467 -17400 -429
rect -17500 -501 -17467 -467
rect -17433 -501 -17400 -467
rect -17500 -539 -17400 -501
rect -17500 -573 -17467 -539
rect -17433 -573 -17400 -539
rect -17500 -611 -17400 -573
rect -17500 -645 -17467 -611
rect -17433 -645 -17400 -611
rect -17500 -683 -17400 -645
rect -17500 -717 -17467 -683
rect -17433 -717 -17400 -683
rect -17500 -755 -17400 -717
rect -17500 -789 -17467 -755
rect -17433 -789 -17400 -755
rect -17500 -827 -17400 -789
rect -17500 -861 -17467 -827
rect -17433 -861 -17400 -827
rect -17500 -899 -17400 -861
rect -17500 -933 -17467 -899
rect -17433 -933 -17400 -899
rect -17500 -971 -17400 -933
rect -17500 -1005 -17467 -971
rect -17433 -1005 -17400 -971
rect -17500 -1043 -17400 -1005
rect -17500 -1077 -17467 -1043
rect -17433 -1077 -17400 -1043
rect -17500 -1115 -17400 -1077
rect -17500 -1149 -17467 -1115
rect -17433 -1149 -17400 -1115
rect -17500 -1187 -17400 -1149
rect -17500 -1221 -17467 -1187
rect -17433 -1221 -17400 -1187
rect -17500 -1259 -17400 -1221
rect -17500 -1293 -17467 -1259
rect -17433 -1293 -17400 -1259
rect -17500 -1331 -17400 -1293
rect -17500 -1365 -17467 -1331
rect -17433 -1365 -17400 -1331
rect -17500 -1403 -17400 -1365
rect -17500 -1437 -17467 -1403
rect -17433 -1437 -17400 -1403
rect -17500 -1475 -17400 -1437
rect -17500 -1509 -17467 -1475
rect -17433 -1509 -17400 -1475
rect -17500 -1547 -17400 -1509
rect -17500 -1581 -17467 -1547
rect -17433 -1581 -17400 -1547
rect -17500 -1619 -17400 -1581
rect -17500 -1653 -17467 -1619
rect -17433 -1653 -17400 -1619
rect -17500 -1691 -17400 -1653
rect -17500 -1725 -17467 -1691
rect -17433 -1725 -17400 -1691
rect -17500 -1763 -17400 -1725
rect -17500 -1797 -17467 -1763
rect -17433 -1780 -17400 -1763
rect 35300 1909 35400 1947
rect 35300 1875 35333 1909
rect 35367 1875 35400 1909
rect 35300 1837 35400 1875
rect 35300 1803 35333 1837
rect 35367 1803 35400 1837
rect 35300 1765 35400 1803
rect 35300 1731 35333 1765
rect 35367 1731 35400 1765
rect 35300 1693 35400 1731
rect 35300 1659 35333 1693
rect 35367 1659 35400 1693
rect 35300 1621 35400 1659
rect 35300 1587 35333 1621
rect 35367 1587 35400 1621
rect 35300 1549 35400 1587
rect 35300 1515 35333 1549
rect 35367 1515 35400 1549
rect 35300 1477 35400 1515
rect 35300 1443 35333 1477
rect 35367 1443 35400 1477
rect 35300 1405 35400 1443
rect 35300 1371 35333 1405
rect 35367 1371 35400 1405
rect 35300 1333 35400 1371
rect 35300 1299 35333 1333
rect 35367 1299 35400 1333
rect 35300 1261 35400 1299
rect 35300 1227 35333 1261
rect 35367 1227 35400 1261
rect 35300 1189 35400 1227
rect 35300 1155 35333 1189
rect 35367 1155 35400 1189
rect 35300 1117 35400 1155
rect 35300 1083 35333 1117
rect 35367 1083 35400 1117
rect 35300 1045 35400 1083
rect 35300 1011 35333 1045
rect 35367 1011 35400 1045
rect 35300 973 35400 1011
rect 35300 939 35333 973
rect 35367 939 35400 973
rect 35300 901 35400 939
rect 35300 867 35333 901
rect 35367 867 35400 901
rect 35300 829 35400 867
rect 35300 795 35333 829
rect 35367 795 35400 829
rect 35300 757 35400 795
rect 35300 723 35333 757
rect 35367 723 35400 757
rect 35300 685 35400 723
rect 35300 651 35333 685
rect 35367 651 35400 685
rect 35300 613 35400 651
rect 35300 579 35333 613
rect 35367 579 35400 613
rect 35300 541 35400 579
rect 35300 507 35333 541
rect 35367 507 35400 541
rect 35300 469 35400 507
rect 35300 435 35333 469
rect 35367 435 35400 469
rect 35300 397 35400 435
rect 35300 363 35333 397
rect 35367 363 35400 397
rect 35300 325 35400 363
rect 35300 291 35333 325
rect 35367 291 35400 325
rect 35300 253 35400 291
rect 35300 219 35333 253
rect 35367 219 35400 253
rect 35300 181 35400 219
rect 35300 147 35333 181
rect 35367 147 35400 181
rect 35300 109 35400 147
rect 35300 75 35333 109
rect 35367 75 35400 109
rect 35300 37 35400 75
rect 35300 3 35333 37
rect 35367 3 35400 37
rect 35300 -35 35400 3
rect 35300 -69 35333 -35
rect 35367 -69 35400 -35
rect 35300 -107 35400 -69
rect 35300 -141 35333 -107
rect 35367 -141 35400 -107
rect 35300 -179 35400 -141
rect 35300 -213 35333 -179
rect 35367 -213 35400 -179
rect 35300 -251 35400 -213
rect 35300 -285 35333 -251
rect 35367 -285 35400 -251
rect 35300 -323 35400 -285
rect 35300 -357 35333 -323
rect 35367 -357 35400 -323
rect 35300 -395 35400 -357
rect 35300 -429 35333 -395
rect 35367 -429 35400 -395
rect 35300 -467 35400 -429
rect 35300 -501 35333 -467
rect 35367 -501 35400 -467
rect 35300 -539 35400 -501
rect 35300 -573 35333 -539
rect 35367 -573 35400 -539
rect 35300 -611 35400 -573
rect 35300 -645 35333 -611
rect 35367 -645 35400 -611
rect 35300 -683 35400 -645
rect 35300 -717 35333 -683
rect 35367 -717 35400 -683
rect 35300 -755 35400 -717
rect 35300 -789 35333 -755
rect 35367 -789 35400 -755
rect 35300 -827 35400 -789
rect 35300 -861 35333 -827
rect 35367 -861 35400 -827
rect 35300 -899 35400 -861
rect 35300 -933 35333 -899
rect 35367 -933 35400 -899
rect 35300 -971 35400 -933
rect 35300 -1005 35333 -971
rect 35367 -1005 35400 -971
rect 35300 -1043 35400 -1005
rect 35300 -1077 35333 -1043
rect 35367 -1077 35400 -1043
rect 35300 -1115 35400 -1077
rect 35300 -1149 35333 -1115
rect 35367 -1149 35400 -1115
rect 35300 -1187 35400 -1149
rect 35300 -1221 35333 -1187
rect 35367 -1221 35400 -1187
rect 35300 -1259 35400 -1221
rect 35300 -1293 35333 -1259
rect 35367 -1293 35400 -1259
rect 35300 -1331 35400 -1293
rect 35300 -1365 35333 -1331
rect 35367 -1365 35400 -1331
rect 35300 -1403 35400 -1365
rect 35300 -1437 35333 -1403
rect 35367 -1437 35400 -1403
rect 35300 -1475 35400 -1437
rect 35300 -1509 35333 -1475
rect 35367 -1509 35400 -1475
rect 35300 -1547 35400 -1509
rect 35300 -1581 35333 -1547
rect 35367 -1581 35400 -1547
rect 35300 -1619 35400 -1581
rect 35300 -1653 35333 -1619
rect 35367 -1653 35400 -1619
rect 35300 -1691 35400 -1653
rect 35300 -1725 35333 -1691
rect 35367 -1725 35400 -1691
rect 35300 -1763 35400 -1725
rect 35300 -1780 35333 -1763
rect -17433 -1797 35333 -1780
rect 35367 -1797 35400 -1763
rect -17500 -1835 35400 -1797
rect -17500 -1869 -17467 -1835
rect -17433 -1860 35333 -1835
rect -17433 -1869 -17400 -1860
rect -17500 -1907 -17400 -1869
rect -17500 -1941 -17467 -1907
rect -17433 -1941 -17400 -1907
rect -17500 -1979 -17400 -1941
rect -17500 -2013 -17467 -1979
rect -17433 -2013 -17400 -1979
rect -17500 -2051 -17400 -2013
rect -17500 -2085 -17467 -2051
rect -17433 -2085 -17400 -2051
rect -17500 -2123 -17400 -2085
rect -17500 -2157 -17467 -2123
rect -17433 -2157 -17400 -2123
rect -17500 -2195 -17400 -2157
rect -17500 -2229 -17467 -2195
rect -17433 -2229 -17400 -2195
rect -17500 -2267 -17400 -2229
rect -17500 -2301 -17467 -2267
rect -17433 -2301 -17400 -2267
rect -17500 -2339 -17400 -2301
rect -17500 -2373 -17467 -2339
rect -17433 -2373 -17400 -2339
rect -17500 -2411 -17400 -2373
rect -17500 -2445 -17467 -2411
rect -17433 -2445 -17400 -2411
rect -17500 -2483 -17400 -2445
rect -17500 -2517 -17467 -2483
rect -17433 -2517 -17400 -2483
rect -17500 -2555 -17400 -2517
rect -17500 -2589 -17467 -2555
rect -17433 -2589 -17400 -2555
rect -17500 -2627 -17400 -2589
rect -17500 -2661 -17467 -2627
rect -17433 -2661 -17400 -2627
rect -17500 -2699 -17400 -2661
rect -17500 -2733 -17467 -2699
rect -17433 -2733 -17400 -2699
rect -17500 -2771 -17400 -2733
rect -17500 -2805 -17467 -2771
rect -17433 -2805 -17400 -2771
rect -17500 -2843 -17400 -2805
rect -17500 -2877 -17467 -2843
rect -17433 -2877 -17400 -2843
rect -17500 -2915 -17400 -2877
rect -17500 -2949 -17467 -2915
rect -17433 -2949 -17400 -2915
rect -17500 -2987 -17400 -2949
rect -17500 -3021 -17467 -2987
rect -17433 -3021 -17400 -2987
rect -17500 -3059 -17400 -3021
rect -17500 -3093 -17467 -3059
rect -17433 -3093 -17400 -3059
rect -17500 -3131 -17400 -3093
rect -17500 -3165 -17467 -3131
rect -17433 -3165 -17400 -3131
rect -17500 -3203 -17400 -3165
rect -17500 -3237 -17467 -3203
rect -17433 -3237 -17400 -3203
rect -17500 -3275 -17400 -3237
rect -17500 -3309 -17467 -3275
rect -17433 -3309 -17400 -3275
rect -17500 -3347 -17400 -3309
rect -17500 -3381 -17467 -3347
rect -17433 -3381 -17400 -3347
rect -17500 -3419 -17400 -3381
rect -17500 -3453 -17467 -3419
rect -17433 -3453 -17400 -3419
rect -17500 -3491 -17400 -3453
rect -17500 -3525 -17467 -3491
rect -17433 -3525 -17400 -3491
rect -17500 -3563 -17400 -3525
rect -17500 -3597 -17467 -3563
rect -17433 -3597 -17400 -3563
rect -17500 -3635 -17400 -3597
rect -17500 -3669 -17467 -3635
rect -17433 -3669 -17400 -3635
rect -17500 -3707 -17400 -3669
rect -17500 -3741 -17467 -3707
rect -17433 -3741 -17400 -3707
rect -17500 -3779 -17400 -3741
rect -17500 -3813 -17467 -3779
rect -17433 -3813 -17400 -3779
rect -17500 -3851 -17400 -3813
rect -17500 -3885 -17467 -3851
rect -17433 -3885 -17400 -3851
rect -17500 -3923 -17400 -3885
rect -17500 -3957 -17467 -3923
rect -17433 -3957 -17400 -3923
rect -17500 -3995 -17400 -3957
rect -17500 -4029 -17467 -3995
rect -17433 -4029 -17400 -3995
rect -17500 -4067 -17400 -4029
rect -17500 -4101 -17467 -4067
rect -17433 -4101 -17400 -4067
rect -17500 -4139 -17400 -4101
rect -17500 -4173 -17467 -4139
rect -17433 -4173 -17400 -4139
rect -17500 -4211 -17400 -4173
rect -17500 -4245 -17467 -4211
rect -17433 -4245 -17400 -4211
rect -17500 -4283 -17400 -4245
rect -17500 -4317 -17467 -4283
rect -17433 -4317 -17400 -4283
rect -17500 -4355 -17400 -4317
rect -17500 -4389 -17467 -4355
rect -17433 -4389 -17400 -4355
rect -17500 -4427 -17400 -4389
rect -17500 -4461 -17467 -4427
rect -17433 -4461 -17400 -4427
rect -17500 -4499 -17400 -4461
rect -17500 -4533 -17467 -4499
rect -17433 -4533 -17400 -4499
rect -17500 -4571 -17400 -4533
rect -17500 -4605 -17467 -4571
rect -17433 -4605 -17400 -4571
rect -17500 -4643 -17400 -4605
rect -17500 -4677 -17467 -4643
rect -17433 -4677 -17400 -4643
rect -17500 -4715 -17400 -4677
rect -17500 -4749 -17467 -4715
rect -17433 -4749 -17400 -4715
rect -17500 -4787 -17400 -4749
rect -17500 -4821 -17467 -4787
rect -17433 -4821 -17400 -4787
rect -17500 -4859 -17400 -4821
rect -17500 -4893 -17467 -4859
rect -17433 -4893 -17400 -4859
rect -17500 -4931 -17400 -4893
rect -17500 -4965 -17467 -4931
rect -17433 -4965 -17400 -4931
rect -17500 -5003 -17400 -4965
rect -17500 -5037 -17467 -5003
rect -17433 -5037 -17400 -5003
rect -17500 -5075 -17400 -5037
rect -17500 -5109 -17467 -5075
rect -17433 -5109 -17400 -5075
rect -17500 -5147 -17400 -5109
rect -17500 -5181 -17467 -5147
rect -17433 -5181 -17400 -5147
rect -17500 -5219 -17400 -5181
rect -17500 -5253 -17467 -5219
rect -17433 -5253 -17400 -5219
rect -17500 -5291 -17400 -5253
rect -17500 -5325 -17467 -5291
rect -17433 -5300 -17400 -5291
rect 35300 -1869 35333 -1860
rect 35367 -1869 35400 -1835
rect 35300 -1907 35400 -1869
rect 35300 -1941 35333 -1907
rect 35367 -1941 35400 -1907
rect 35300 -1979 35400 -1941
rect 35300 -2013 35333 -1979
rect 35367 -2013 35400 -1979
rect 35300 -2051 35400 -2013
rect 35300 -2085 35333 -2051
rect 35367 -2085 35400 -2051
rect 35300 -2123 35400 -2085
rect 35300 -2157 35333 -2123
rect 35367 -2157 35400 -2123
rect 35300 -2195 35400 -2157
rect 35300 -2229 35333 -2195
rect 35367 -2229 35400 -2195
rect 35300 -2267 35400 -2229
rect 35300 -2301 35333 -2267
rect 35367 -2301 35400 -2267
rect 35300 -2339 35400 -2301
rect 35300 -2373 35333 -2339
rect 35367 -2373 35400 -2339
rect 35300 -2411 35400 -2373
rect 35300 -2445 35333 -2411
rect 35367 -2445 35400 -2411
rect 35300 -2483 35400 -2445
rect 35300 -2517 35333 -2483
rect 35367 -2517 35400 -2483
rect 35300 -2555 35400 -2517
rect 35300 -2589 35333 -2555
rect 35367 -2589 35400 -2555
rect 35300 -2627 35400 -2589
rect 35300 -2661 35333 -2627
rect 35367 -2661 35400 -2627
rect 35300 -2699 35400 -2661
rect 35300 -2733 35333 -2699
rect 35367 -2733 35400 -2699
rect 35300 -2771 35400 -2733
rect 35300 -2805 35333 -2771
rect 35367 -2805 35400 -2771
rect 35300 -2843 35400 -2805
rect 35300 -2877 35333 -2843
rect 35367 -2877 35400 -2843
rect 35300 -2915 35400 -2877
rect 35300 -2949 35333 -2915
rect 35367 -2949 35400 -2915
rect 35300 -2987 35400 -2949
rect 35300 -3021 35333 -2987
rect 35367 -3021 35400 -2987
rect 35300 -3059 35400 -3021
rect 35300 -3093 35333 -3059
rect 35367 -3093 35400 -3059
rect 35300 -3131 35400 -3093
rect 35300 -3165 35333 -3131
rect 35367 -3165 35400 -3131
rect 35300 -3203 35400 -3165
rect 35300 -3237 35333 -3203
rect 35367 -3237 35400 -3203
rect 35300 -3275 35400 -3237
rect 35300 -3309 35333 -3275
rect 35367 -3309 35400 -3275
rect 35300 -3347 35400 -3309
rect 35300 -3381 35333 -3347
rect 35367 -3381 35400 -3347
rect 35300 -3419 35400 -3381
rect 35300 -3453 35333 -3419
rect 35367 -3453 35400 -3419
rect 35300 -3491 35400 -3453
rect 35300 -3525 35333 -3491
rect 35367 -3525 35400 -3491
rect 35300 -3563 35400 -3525
rect 35300 -3597 35333 -3563
rect 35367 -3597 35400 -3563
rect 35300 -3635 35400 -3597
rect 35300 -3669 35333 -3635
rect 35367 -3669 35400 -3635
rect 35300 -3707 35400 -3669
rect 35300 -3741 35333 -3707
rect 35367 -3741 35400 -3707
rect 35300 -3779 35400 -3741
rect 35300 -3813 35333 -3779
rect 35367 -3813 35400 -3779
rect 35300 -3851 35400 -3813
rect 35300 -3885 35333 -3851
rect 35367 -3885 35400 -3851
rect 35300 -3923 35400 -3885
rect 35300 -3957 35333 -3923
rect 35367 -3957 35400 -3923
rect 35300 -3995 35400 -3957
rect 35300 -4029 35333 -3995
rect 35367 -4029 35400 -3995
rect 35300 -4067 35400 -4029
rect 35300 -4101 35333 -4067
rect 35367 -4101 35400 -4067
rect 35300 -4139 35400 -4101
rect 35300 -4173 35333 -4139
rect 35367 -4173 35400 -4139
rect 35300 -4211 35400 -4173
rect 35300 -4245 35333 -4211
rect 35367 -4245 35400 -4211
rect 35300 -4283 35400 -4245
rect 35300 -4317 35333 -4283
rect 35367 -4317 35400 -4283
rect 35300 -4355 35400 -4317
rect 35300 -4389 35333 -4355
rect 35367 -4389 35400 -4355
rect 35300 -4427 35400 -4389
rect 35300 -4461 35333 -4427
rect 35367 -4461 35400 -4427
rect 35300 -4499 35400 -4461
rect 35300 -4533 35333 -4499
rect 35367 -4533 35400 -4499
rect 35300 -4571 35400 -4533
rect 35300 -4605 35333 -4571
rect 35367 -4605 35400 -4571
rect 35300 -4643 35400 -4605
rect 35300 -4677 35333 -4643
rect 35367 -4677 35400 -4643
rect 35300 -4715 35400 -4677
rect 35300 -4749 35333 -4715
rect 35367 -4749 35400 -4715
rect 35300 -4787 35400 -4749
rect 35300 -4821 35333 -4787
rect 35367 -4821 35400 -4787
rect 35300 -4859 35400 -4821
rect 35300 -4893 35333 -4859
rect 35367 -4893 35400 -4859
rect 35300 -4931 35400 -4893
rect 35300 -4965 35333 -4931
rect 35367 -4965 35400 -4931
rect 35300 -5003 35400 -4965
rect 35300 -5037 35333 -5003
rect 35367 -5037 35400 -5003
rect 35300 -5075 35400 -5037
rect 35300 -5109 35333 -5075
rect 35367 -5109 35400 -5075
rect 35300 -5147 35400 -5109
rect 35300 -5181 35333 -5147
rect 35367 -5181 35400 -5147
rect 35300 -5219 35400 -5181
rect 35300 -5253 35333 -5219
rect 35367 -5253 35400 -5219
rect 35300 -5291 35400 -5253
rect 35300 -5300 35333 -5291
rect -17433 -5325 35333 -5300
rect 35367 -5325 35400 -5291
rect -17500 -5363 35400 -5325
rect -17500 -5397 -17467 -5363
rect -17433 -5380 35333 -5363
rect -17433 -5397 -17400 -5380
rect -17500 -5435 -17400 -5397
rect -17500 -5469 -17467 -5435
rect -17433 -5469 -17400 -5435
rect -17500 -5507 -17400 -5469
rect -17500 -5541 -17467 -5507
rect -17433 -5541 -17400 -5507
rect -17500 -5579 -17400 -5541
rect -17500 -5613 -17467 -5579
rect -17433 -5613 -17400 -5579
rect -17500 -5651 -17400 -5613
rect -17500 -5685 -17467 -5651
rect -17433 -5685 -17400 -5651
rect -17500 -5723 -17400 -5685
rect -17500 -5757 -17467 -5723
rect -17433 -5757 -17400 -5723
rect -17500 -5795 -17400 -5757
rect -17500 -5829 -17467 -5795
rect -17433 -5829 -17400 -5795
rect -17500 -5867 -17400 -5829
rect -17500 -5901 -17467 -5867
rect -17433 -5901 -17400 -5867
rect -17500 -5939 -17400 -5901
rect -17500 -5973 -17467 -5939
rect -17433 -5973 -17400 -5939
rect -17500 -6011 -17400 -5973
rect -17500 -6045 -17467 -6011
rect -17433 -6045 -17400 -6011
rect -17500 -6083 -17400 -6045
rect -17500 -6117 -17467 -6083
rect -17433 -6117 -17400 -6083
rect -17500 -6155 -17400 -6117
rect -17500 -6189 -17467 -6155
rect -17433 -6189 -17400 -6155
rect -17500 -6227 -17400 -6189
rect -17500 -6261 -17467 -6227
rect -17433 -6261 -17400 -6227
rect -17500 -6299 -17400 -6261
rect -17500 -6333 -17467 -6299
rect -17433 -6333 -17400 -6299
rect -17500 -6371 -17400 -6333
rect -17500 -6405 -17467 -6371
rect -17433 -6405 -17400 -6371
rect -17500 -6443 -17400 -6405
rect -17500 -6477 -17467 -6443
rect -17433 -6477 -17400 -6443
rect -17500 -6515 -17400 -6477
rect -17500 -6549 -17467 -6515
rect -17433 -6549 -17400 -6515
rect -17500 -6587 -17400 -6549
rect -17500 -6621 -17467 -6587
rect -17433 -6621 -17400 -6587
rect -17500 -6659 -17400 -6621
rect -17500 -6693 -17467 -6659
rect -17433 -6693 -17400 -6659
rect -17500 -6731 -17400 -6693
rect -17500 -6765 -17467 -6731
rect -17433 -6765 -17400 -6731
rect -17500 -6803 -17400 -6765
rect -17500 -6837 -17467 -6803
rect -17433 -6837 -17400 -6803
rect -17500 -6875 -17400 -6837
rect -17500 -6909 -17467 -6875
rect -17433 -6909 -17400 -6875
rect -17500 -6947 -17400 -6909
rect -17500 -6981 -17467 -6947
rect -17433 -6981 -17400 -6947
rect -17500 -7019 -17400 -6981
rect -17500 -7053 -17467 -7019
rect -17433 -7053 -17400 -7019
rect -17500 -7091 -17400 -7053
rect -17500 -7125 -17467 -7091
rect -17433 -7125 -17400 -7091
rect -17500 -7163 -17400 -7125
rect -17500 -7197 -17467 -7163
rect -17433 -7197 -17400 -7163
rect -17500 -7200 -17400 -7197
rect 35300 -5397 35333 -5380
rect 35367 -5397 35400 -5363
rect 35300 -5435 35400 -5397
rect 35300 -5469 35333 -5435
rect 35367 -5469 35400 -5435
rect 35300 -5507 35400 -5469
rect 35300 -5541 35333 -5507
rect 35367 -5541 35400 -5507
rect 35300 -5579 35400 -5541
rect 35300 -5613 35333 -5579
rect 35367 -5613 35400 -5579
rect 35300 -5651 35400 -5613
rect 35300 -5685 35333 -5651
rect 35367 -5685 35400 -5651
rect 35300 -5723 35400 -5685
rect 35300 -5757 35333 -5723
rect 35367 -5757 35400 -5723
rect 35300 -5795 35400 -5757
rect 35300 -5829 35333 -5795
rect 35367 -5829 35400 -5795
rect 35300 -5867 35400 -5829
rect 35300 -5901 35333 -5867
rect 35367 -5901 35400 -5867
rect 35300 -5939 35400 -5901
rect 35300 -5973 35333 -5939
rect 35367 -5973 35400 -5939
rect 35300 -6011 35400 -5973
rect 35300 -6045 35333 -6011
rect 35367 -6045 35400 -6011
rect 35300 -6083 35400 -6045
rect 35300 -6117 35333 -6083
rect 35367 -6117 35400 -6083
rect 35300 -6155 35400 -6117
rect 35300 -6189 35333 -6155
rect 35367 -6189 35400 -6155
rect 35300 -6227 35400 -6189
rect 35300 -6261 35333 -6227
rect 35367 -6261 35400 -6227
rect 35300 -6299 35400 -6261
rect 35300 -6333 35333 -6299
rect 35367 -6333 35400 -6299
rect 35300 -6371 35400 -6333
rect 35300 -6405 35333 -6371
rect 35367 -6405 35400 -6371
rect 35300 -6443 35400 -6405
rect 35300 -6477 35333 -6443
rect 35367 -6477 35400 -6443
rect 35300 -6515 35400 -6477
rect 35300 -6549 35333 -6515
rect 35367 -6549 35400 -6515
rect 35300 -6587 35400 -6549
rect 35300 -6621 35333 -6587
rect 35367 -6621 35400 -6587
rect 35300 -6659 35400 -6621
rect 35300 -6693 35333 -6659
rect 35367 -6693 35400 -6659
rect 35300 -6731 35400 -6693
rect 35300 -6765 35333 -6731
rect 35367 -6765 35400 -6731
rect 35300 -6803 35400 -6765
rect 35300 -6837 35333 -6803
rect 35367 -6837 35400 -6803
rect 35300 -6875 35400 -6837
rect 35300 -6909 35333 -6875
rect 35367 -6909 35400 -6875
rect 35300 -6947 35400 -6909
rect 35300 -6981 35333 -6947
rect 35367 -6981 35400 -6947
rect 35300 -7019 35400 -6981
rect 35300 -7053 35333 -7019
rect 35367 -7053 35400 -7019
rect 35300 -7091 35400 -7053
rect 35300 -7125 35333 -7091
rect 35367 -7125 35400 -7091
rect 35300 -7163 35400 -7125
rect 35300 -7197 35333 -7163
rect 35367 -7197 35400 -7163
rect 35300 -7200 35400 -7197
rect -17500 -7233 35400 -7200
rect -17500 -7267 -17321 -7233
rect -17287 -7267 -17249 -7233
rect -17215 -7267 -17177 -7233
rect -17143 -7267 -17105 -7233
rect -17071 -7267 -17033 -7233
rect -16999 -7267 -16961 -7233
rect -16927 -7267 -16889 -7233
rect -16855 -7267 -16817 -7233
rect -16783 -7267 -16745 -7233
rect -16711 -7267 -16673 -7233
rect -16639 -7267 -16601 -7233
rect -16567 -7267 -16529 -7233
rect -16495 -7267 -16457 -7233
rect -16423 -7267 -16385 -7233
rect -16351 -7267 -16313 -7233
rect -16279 -7267 -16241 -7233
rect -16207 -7267 -16169 -7233
rect -16135 -7267 -16097 -7233
rect -16063 -7267 -16025 -7233
rect -15991 -7267 -15953 -7233
rect -15919 -7267 -15881 -7233
rect -15847 -7267 -15809 -7233
rect -15775 -7267 -15737 -7233
rect -15703 -7267 -15665 -7233
rect -15631 -7267 -15593 -7233
rect -15559 -7267 -15521 -7233
rect -15487 -7267 -15449 -7233
rect -15415 -7267 -15377 -7233
rect -15343 -7267 -15305 -7233
rect -15271 -7267 -15233 -7233
rect -15199 -7267 -15161 -7233
rect -15127 -7267 -15089 -7233
rect -15055 -7267 -15017 -7233
rect -14983 -7267 -14945 -7233
rect -14911 -7267 -14873 -7233
rect -14839 -7267 -14801 -7233
rect -14767 -7267 -14729 -7233
rect -14695 -7267 -14657 -7233
rect -14623 -7267 -14585 -7233
rect -14551 -7267 -14513 -7233
rect -14479 -7267 -14441 -7233
rect -14407 -7267 -14369 -7233
rect -14335 -7267 -14297 -7233
rect -14263 -7267 -14225 -7233
rect -14191 -7267 -14153 -7233
rect -14119 -7267 -14081 -7233
rect -14047 -7267 -14009 -7233
rect -13975 -7267 -13937 -7233
rect -13903 -7267 -13865 -7233
rect -13831 -7267 -13793 -7233
rect -13759 -7267 -13721 -7233
rect -13687 -7267 -13649 -7233
rect -13615 -7267 -13577 -7233
rect -13543 -7267 -13505 -7233
rect -13471 -7267 -13433 -7233
rect -13399 -7267 -13361 -7233
rect -13327 -7267 -13289 -7233
rect -13255 -7267 -13217 -7233
rect -13183 -7267 -13145 -7233
rect -13111 -7267 -13073 -7233
rect -13039 -7267 -13001 -7233
rect -12967 -7267 -12929 -7233
rect -12895 -7267 -12857 -7233
rect -12823 -7267 -12785 -7233
rect -12751 -7267 -12713 -7233
rect -12679 -7267 -12641 -7233
rect -12607 -7267 -12569 -7233
rect -12535 -7267 -12497 -7233
rect -12463 -7267 -12425 -7233
rect -12391 -7267 -12353 -7233
rect -12319 -7267 -12281 -7233
rect -12247 -7267 -12209 -7233
rect -12175 -7267 -12137 -7233
rect -12103 -7267 -12065 -7233
rect -12031 -7267 -11993 -7233
rect -11959 -7267 -11921 -7233
rect -11887 -7267 -11849 -7233
rect -11815 -7267 -11777 -7233
rect -11743 -7267 -11705 -7233
rect -11671 -7267 -11633 -7233
rect -11599 -7267 -11561 -7233
rect -11527 -7267 -11489 -7233
rect -11455 -7267 -11417 -7233
rect -11383 -7267 -11345 -7233
rect -11311 -7267 -11273 -7233
rect -11239 -7267 -11201 -7233
rect -11167 -7267 -11129 -7233
rect -11095 -7267 -11057 -7233
rect -11023 -7267 -10985 -7233
rect -10951 -7267 -10913 -7233
rect -10879 -7267 -10841 -7233
rect -10807 -7267 -10769 -7233
rect -10735 -7267 -10697 -7233
rect -10663 -7267 -10625 -7233
rect -10591 -7267 -10553 -7233
rect -10519 -7267 -10481 -7233
rect -10447 -7267 -10409 -7233
rect -10375 -7267 -10337 -7233
rect -10303 -7267 -10265 -7233
rect -10231 -7267 -10193 -7233
rect -10159 -7267 -10121 -7233
rect -10087 -7267 -10049 -7233
rect -10015 -7267 -9977 -7233
rect -9943 -7267 -9905 -7233
rect -9871 -7267 -9833 -7233
rect -9799 -7267 -9761 -7233
rect -9727 -7267 -9689 -7233
rect -9655 -7267 -9617 -7233
rect -9583 -7267 -9545 -7233
rect -9511 -7267 -9473 -7233
rect -9439 -7267 -9401 -7233
rect -9367 -7267 -9329 -7233
rect -9295 -7267 -9257 -7233
rect -9223 -7267 -9185 -7233
rect -9151 -7267 -9113 -7233
rect -9079 -7267 -9041 -7233
rect -9007 -7267 -8969 -7233
rect -8935 -7267 -8897 -7233
rect -8863 -7267 -8825 -7233
rect -8791 -7267 -8753 -7233
rect -8719 -7267 -8681 -7233
rect -8647 -7267 -8609 -7233
rect -8575 -7267 -8537 -7233
rect -8503 -7267 -8465 -7233
rect -8431 -7267 -8393 -7233
rect -8359 -7267 -8321 -7233
rect -8287 -7267 -8249 -7233
rect -8215 -7267 -8177 -7233
rect -8143 -7267 -8105 -7233
rect -8071 -7267 -8033 -7233
rect -7999 -7267 -7961 -7233
rect -7927 -7267 -7889 -7233
rect -7855 -7267 -7817 -7233
rect -7783 -7267 -7745 -7233
rect -7711 -7267 -7673 -7233
rect -7639 -7267 -7601 -7233
rect -7567 -7267 -7529 -7233
rect -7495 -7267 -7457 -7233
rect -7423 -7267 -7385 -7233
rect -7351 -7267 -7313 -7233
rect -7279 -7267 -7241 -7233
rect -7207 -7267 -7169 -7233
rect -7135 -7267 -7097 -7233
rect -7063 -7267 -7025 -7233
rect -6991 -7267 -6953 -7233
rect -6919 -7267 -6881 -7233
rect -6847 -7267 -6809 -7233
rect -6775 -7267 -6737 -7233
rect -6703 -7267 -6665 -7233
rect -6631 -7267 -6593 -7233
rect -6559 -7267 -6521 -7233
rect -6487 -7267 -6449 -7233
rect -6415 -7267 -6377 -7233
rect -6343 -7267 -6305 -7233
rect -6271 -7267 -6233 -7233
rect -6199 -7267 -6161 -7233
rect -6127 -7267 -6089 -7233
rect -6055 -7267 -6017 -7233
rect -5983 -7267 -5945 -7233
rect -5911 -7267 -5873 -7233
rect -5839 -7267 -5801 -7233
rect -5767 -7267 -5729 -7233
rect -5695 -7267 -5657 -7233
rect -5623 -7267 -5585 -7233
rect -5551 -7267 -5513 -7233
rect -5479 -7267 -5441 -7233
rect -5407 -7267 -5369 -7233
rect -5335 -7267 -5297 -7233
rect -5263 -7267 -5225 -7233
rect -5191 -7267 -5153 -7233
rect -5119 -7267 -5081 -7233
rect -5047 -7267 -5009 -7233
rect -4975 -7267 -4937 -7233
rect -4903 -7267 -4865 -7233
rect -4831 -7267 -4793 -7233
rect -4759 -7267 -4721 -7233
rect -4687 -7267 -4649 -7233
rect -4615 -7267 -4577 -7233
rect -4543 -7267 -4505 -7233
rect -4471 -7267 -4433 -7233
rect -4399 -7267 -4361 -7233
rect -4327 -7267 -4289 -7233
rect -4255 -7267 -4217 -7233
rect -4183 -7267 -4145 -7233
rect -4111 -7267 -4073 -7233
rect -4039 -7267 -4001 -7233
rect -3967 -7267 -3929 -7233
rect -3895 -7267 -3857 -7233
rect -3823 -7267 -3785 -7233
rect -3751 -7267 -3713 -7233
rect -3679 -7267 -3641 -7233
rect -3607 -7267 -3569 -7233
rect -3535 -7267 -3497 -7233
rect -3463 -7267 -3425 -7233
rect -3391 -7267 -3353 -7233
rect -3319 -7267 -3281 -7233
rect -3247 -7267 -3209 -7233
rect -3175 -7267 -3137 -7233
rect -3103 -7267 -3065 -7233
rect -3031 -7267 -2993 -7233
rect -2959 -7267 -2921 -7233
rect -2887 -7267 -2849 -7233
rect -2815 -7267 -2777 -7233
rect -2743 -7267 -2705 -7233
rect -2671 -7267 -2633 -7233
rect -2599 -7267 -2561 -7233
rect -2527 -7267 -2489 -7233
rect -2455 -7267 -2417 -7233
rect -2383 -7267 -2345 -7233
rect -2311 -7267 -2273 -7233
rect -2239 -7267 -2201 -7233
rect -2167 -7267 -2129 -7233
rect -2095 -7267 -2057 -7233
rect -2023 -7267 -1985 -7233
rect -1951 -7267 -1913 -7233
rect -1879 -7267 -1841 -7233
rect -1807 -7267 -1769 -7233
rect -1735 -7267 -1697 -7233
rect -1663 -7267 -1625 -7233
rect -1591 -7267 -1553 -7233
rect -1519 -7267 -1481 -7233
rect -1447 -7267 -1409 -7233
rect -1375 -7267 -1337 -7233
rect -1303 -7267 -1265 -7233
rect -1231 -7267 -1193 -7233
rect -1159 -7267 -1121 -7233
rect -1087 -7267 -1049 -7233
rect -1015 -7267 -977 -7233
rect -943 -7267 -905 -7233
rect -871 -7267 -833 -7233
rect -799 -7267 -761 -7233
rect -727 -7267 -689 -7233
rect -655 -7267 -617 -7233
rect -583 -7267 -545 -7233
rect -511 -7267 -473 -7233
rect -439 -7267 -401 -7233
rect -367 -7267 -329 -7233
rect -295 -7267 -257 -7233
rect -223 -7267 -185 -7233
rect -151 -7267 -113 -7233
rect -79 -7267 -41 -7233
rect -7 -7267 31 -7233
rect 65 -7267 103 -7233
rect 137 -7267 175 -7233
rect 209 -7267 247 -7233
rect 281 -7267 319 -7233
rect 353 -7267 391 -7233
rect 425 -7267 463 -7233
rect 497 -7267 535 -7233
rect 569 -7267 607 -7233
rect 641 -7267 679 -7233
rect 713 -7267 751 -7233
rect 785 -7267 823 -7233
rect 857 -7267 895 -7233
rect 929 -7267 967 -7233
rect 1001 -7267 1039 -7233
rect 1073 -7267 1111 -7233
rect 1145 -7267 1183 -7233
rect 1217 -7267 1255 -7233
rect 1289 -7267 1327 -7233
rect 1361 -7267 1399 -7233
rect 1433 -7267 1471 -7233
rect 1505 -7267 1543 -7233
rect 1577 -7267 1615 -7233
rect 1649 -7267 1687 -7233
rect 1721 -7267 1759 -7233
rect 1793 -7267 1831 -7233
rect 1865 -7267 1903 -7233
rect 1937 -7267 1975 -7233
rect 2009 -7267 2047 -7233
rect 2081 -7267 2119 -7233
rect 2153 -7267 2191 -7233
rect 2225 -7267 2263 -7233
rect 2297 -7267 2335 -7233
rect 2369 -7267 2407 -7233
rect 2441 -7267 2479 -7233
rect 2513 -7267 2551 -7233
rect 2585 -7267 2623 -7233
rect 2657 -7267 2695 -7233
rect 2729 -7267 2767 -7233
rect 2801 -7267 2839 -7233
rect 2873 -7267 2911 -7233
rect 2945 -7267 2983 -7233
rect 3017 -7267 3055 -7233
rect 3089 -7267 3127 -7233
rect 3161 -7267 3199 -7233
rect 3233 -7267 3271 -7233
rect 3305 -7267 3343 -7233
rect 3377 -7267 3415 -7233
rect 3449 -7267 3487 -7233
rect 3521 -7267 3559 -7233
rect 3593 -7267 3631 -7233
rect 3665 -7267 3703 -7233
rect 3737 -7267 3775 -7233
rect 3809 -7267 3847 -7233
rect 3881 -7267 3919 -7233
rect 3953 -7267 3991 -7233
rect 4025 -7267 4063 -7233
rect 4097 -7267 4135 -7233
rect 4169 -7267 4207 -7233
rect 4241 -7267 4279 -7233
rect 4313 -7267 4351 -7233
rect 4385 -7267 4423 -7233
rect 4457 -7267 4495 -7233
rect 4529 -7267 4567 -7233
rect 4601 -7267 4639 -7233
rect 4673 -7267 4711 -7233
rect 4745 -7267 4783 -7233
rect 4817 -7267 4855 -7233
rect 4889 -7267 4927 -7233
rect 4961 -7267 4999 -7233
rect 5033 -7267 5071 -7233
rect 5105 -7267 5143 -7233
rect 5177 -7267 5215 -7233
rect 5249 -7267 5287 -7233
rect 5321 -7267 5359 -7233
rect 5393 -7267 5431 -7233
rect 5465 -7267 5503 -7233
rect 5537 -7267 5575 -7233
rect 5609 -7267 5647 -7233
rect 5681 -7267 5719 -7233
rect 5753 -7267 5791 -7233
rect 5825 -7267 5863 -7233
rect 5897 -7267 5935 -7233
rect 5969 -7267 6007 -7233
rect 6041 -7267 6079 -7233
rect 6113 -7267 6151 -7233
rect 6185 -7267 6223 -7233
rect 6257 -7267 6295 -7233
rect 6329 -7267 6367 -7233
rect 6401 -7267 6439 -7233
rect 6473 -7267 6511 -7233
rect 6545 -7267 6583 -7233
rect 6617 -7267 6655 -7233
rect 6689 -7267 6727 -7233
rect 6761 -7267 6799 -7233
rect 6833 -7267 6871 -7233
rect 6905 -7267 6943 -7233
rect 6977 -7267 7015 -7233
rect 7049 -7267 7087 -7233
rect 7121 -7267 7159 -7233
rect 7193 -7267 7231 -7233
rect 7265 -7267 7303 -7233
rect 7337 -7267 7375 -7233
rect 7409 -7267 7447 -7233
rect 7481 -7267 7519 -7233
rect 7553 -7267 7591 -7233
rect 7625 -7267 7663 -7233
rect 7697 -7267 7735 -7233
rect 7769 -7267 7807 -7233
rect 7841 -7267 7879 -7233
rect 7913 -7267 7951 -7233
rect 7985 -7267 8023 -7233
rect 8057 -7267 8095 -7233
rect 8129 -7267 8167 -7233
rect 8201 -7267 8239 -7233
rect 8273 -7267 8311 -7233
rect 8345 -7267 8383 -7233
rect 8417 -7267 8455 -7233
rect 8489 -7267 8527 -7233
rect 8561 -7267 8599 -7233
rect 8633 -7267 8671 -7233
rect 8705 -7267 8743 -7233
rect 8777 -7267 8815 -7233
rect 8849 -7267 8887 -7233
rect 8921 -7267 8959 -7233
rect 8993 -7267 9031 -7233
rect 9065 -7267 9103 -7233
rect 9137 -7267 9175 -7233
rect 9209 -7267 9247 -7233
rect 9281 -7267 9319 -7233
rect 9353 -7267 9391 -7233
rect 9425 -7267 9463 -7233
rect 9497 -7267 9535 -7233
rect 9569 -7267 9607 -7233
rect 9641 -7267 9679 -7233
rect 9713 -7267 9751 -7233
rect 9785 -7267 9823 -7233
rect 9857 -7267 9895 -7233
rect 9929 -7267 9967 -7233
rect 10001 -7267 10039 -7233
rect 10073 -7267 10111 -7233
rect 10145 -7267 10183 -7233
rect 10217 -7267 10255 -7233
rect 10289 -7267 10327 -7233
rect 10361 -7267 10399 -7233
rect 10433 -7267 10471 -7233
rect 10505 -7267 10543 -7233
rect 10577 -7267 10615 -7233
rect 10649 -7267 10687 -7233
rect 10721 -7267 10759 -7233
rect 10793 -7267 10831 -7233
rect 10865 -7267 10903 -7233
rect 10937 -7267 10975 -7233
rect 11009 -7267 11047 -7233
rect 11081 -7267 11119 -7233
rect 11153 -7267 11191 -7233
rect 11225 -7267 11263 -7233
rect 11297 -7267 11335 -7233
rect 11369 -7267 11407 -7233
rect 11441 -7267 11479 -7233
rect 11513 -7267 11551 -7233
rect 11585 -7267 11623 -7233
rect 11657 -7267 11695 -7233
rect 11729 -7267 11767 -7233
rect 11801 -7267 11839 -7233
rect 11873 -7267 11911 -7233
rect 11945 -7267 11983 -7233
rect 12017 -7267 12055 -7233
rect 12089 -7267 12127 -7233
rect 12161 -7267 12199 -7233
rect 12233 -7267 12271 -7233
rect 12305 -7267 12343 -7233
rect 12377 -7267 12415 -7233
rect 12449 -7267 12487 -7233
rect 12521 -7267 12559 -7233
rect 12593 -7267 12631 -7233
rect 12665 -7267 12703 -7233
rect 12737 -7267 12775 -7233
rect 12809 -7267 12847 -7233
rect 12881 -7267 12919 -7233
rect 12953 -7267 12991 -7233
rect 13025 -7267 13063 -7233
rect 13097 -7267 13135 -7233
rect 13169 -7267 13207 -7233
rect 13241 -7267 13279 -7233
rect 13313 -7267 13351 -7233
rect 13385 -7267 13423 -7233
rect 13457 -7267 13495 -7233
rect 13529 -7267 13567 -7233
rect 13601 -7267 13639 -7233
rect 13673 -7267 13711 -7233
rect 13745 -7267 13783 -7233
rect 13817 -7267 13855 -7233
rect 13889 -7267 13927 -7233
rect 13961 -7267 13999 -7233
rect 14033 -7267 14071 -7233
rect 14105 -7267 14143 -7233
rect 14177 -7267 14215 -7233
rect 14249 -7267 14287 -7233
rect 14321 -7267 14359 -7233
rect 14393 -7267 14431 -7233
rect 14465 -7267 14503 -7233
rect 14537 -7267 14575 -7233
rect 14609 -7267 14647 -7233
rect 14681 -7267 14719 -7233
rect 14753 -7267 14791 -7233
rect 14825 -7267 14863 -7233
rect 14897 -7267 14935 -7233
rect 14969 -7267 15007 -7233
rect 15041 -7267 15079 -7233
rect 15113 -7267 15151 -7233
rect 15185 -7267 15223 -7233
rect 15257 -7267 15295 -7233
rect 15329 -7267 15367 -7233
rect 15401 -7267 15439 -7233
rect 15473 -7267 15511 -7233
rect 15545 -7267 15583 -7233
rect 15617 -7267 15655 -7233
rect 15689 -7267 15727 -7233
rect 15761 -7267 15799 -7233
rect 15833 -7267 15871 -7233
rect 15905 -7267 15943 -7233
rect 15977 -7267 16015 -7233
rect 16049 -7267 16087 -7233
rect 16121 -7267 16159 -7233
rect 16193 -7267 16231 -7233
rect 16265 -7267 16303 -7233
rect 16337 -7267 16375 -7233
rect 16409 -7267 16447 -7233
rect 16481 -7267 16519 -7233
rect 16553 -7267 16591 -7233
rect 16625 -7267 16663 -7233
rect 16697 -7267 16735 -7233
rect 16769 -7267 16807 -7233
rect 16841 -7267 16879 -7233
rect 16913 -7267 16951 -7233
rect 16985 -7267 17023 -7233
rect 17057 -7267 17095 -7233
rect 17129 -7267 17167 -7233
rect 17201 -7267 17239 -7233
rect 17273 -7267 17311 -7233
rect 17345 -7267 17383 -7233
rect 17417 -7267 17455 -7233
rect 17489 -7267 17527 -7233
rect 17561 -7267 17599 -7233
rect 17633 -7267 17671 -7233
rect 17705 -7267 17743 -7233
rect 17777 -7267 17815 -7233
rect 17849 -7267 17887 -7233
rect 17921 -7267 17959 -7233
rect 17993 -7267 18031 -7233
rect 18065 -7267 18103 -7233
rect 18137 -7267 18175 -7233
rect 18209 -7267 18247 -7233
rect 18281 -7267 18319 -7233
rect 18353 -7267 18391 -7233
rect 18425 -7267 18463 -7233
rect 18497 -7267 18535 -7233
rect 18569 -7267 18607 -7233
rect 18641 -7267 18679 -7233
rect 18713 -7267 18751 -7233
rect 18785 -7267 18823 -7233
rect 18857 -7267 18895 -7233
rect 18929 -7267 18967 -7233
rect 19001 -7267 19039 -7233
rect 19073 -7267 19111 -7233
rect 19145 -7267 19183 -7233
rect 19217 -7267 19255 -7233
rect 19289 -7267 19327 -7233
rect 19361 -7267 19399 -7233
rect 19433 -7267 19471 -7233
rect 19505 -7267 19543 -7233
rect 19577 -7267 19615 -7233
rect 19649 -7267 19687 -7233
rect 19721 -7267 19759 -7233
rect 19793 -7267 19831 -7233
rect 19865 -7267 19903 -7233
rect 19937 -7267 19975 -7233
rect 20009 -7267 20047 -7233
rect 20081 -7267 20119 -7233
rect 20153 -7267 20191 -7233
rect 20225 -7267 20263 -7233
rect 20297 -7267 20335 -7233
rect 20369 -7267 20407 -7233
rect 20441 -7267 20479 -7233
rect 20513 -7267 20551 -7233
rect 20585 -7267 20623 -7233
rect 20657 -7267 20695 -7233
rect 20729 -7267 20767 -7233
rect 20801 -7267 20839 -7233
rect 20873 -7267 20911 -7233
rect 20945 -7267 20983 -7233
rect 21017 -7267 21055 -7233
rect 21089 -7267 21127 -7233
rect 21161 -7267 21199 -7233
rect 21233 -7267 21271 -7233
rect 21305 -7267 21343 -7233
rect 21377 -7267 21415 -7233
rect 21449 -7267 21487 -7233
rect 21521 -7267 21559 -7233
rect 21593 -7267 21631 -7233
rect 21665 -7267 21703 -7233
rect 21737 -7267 21775 -7233
rect 21809 -7267 21847 -7233
rect 21881 -7267 21919 -7233
rect 21953 -7267 21991 -7233
rect 22025 -7267 22063 -7233
rect 22097 -7267 22135 -7233
rect 22169 -7267 22207 -7233
rect 22241 -7267 22279 -7233
rect 22313 -7267 22351 -7233
rect 22385 -7267 22423 -7233
rect 22457 -7267 22495 -7233
rect 22529 -7267 22567 -7233
rect 22601 -7267 22639 -7233
rect 22673 -7267 22711 -7233
rect 22745 -7267 22783 -7233
rect 22817 -7267 22855 -7233
rect 22889 -7267 22927 -7233
rect 22961 -7267 22999 -7233
rect 23033 -7267 23071 -7233
rect 23105 -7267 23143 -7233
rect 23177 -7267 23215 -7233
rect 23249 -7267 23287 -7233
rect 23321 -7267 23359 -7233
rect 23393 -7267 23431 -7233
rect 23465 -7267 23503 -7233
rect 23537 -7267 23575 -7233
rect 23609 -7267 23647 -7233
rect 23681 -7267 23719 -7233
rect 23753 -7267 23791 -7233
rect 23825 -7267 23863 -7233
rect 23897 -7267 23935 -7233
rect 23969 -7267 24007 -7233
rect 24041 -7267 24079 -7233
rect 24113 -7267 24151 -7233
rect 24185 -7267 24223 -7233
rect 24257 -7267 24295 -7233
rect 24329 -7267 24367 -7233
rect 24401 -7267 24439 -7233
rect 24473 -7267 24511 -7233
rect 24545 -7267 24583 -7233
rect 24617 -7267 24655 -7233
rect 24689 -7267 24727 -7233
rect 24761 -7267 24799 -7233
rect 24833 -7267 24871 -7233
rect 24905 -7267 24943 -7233
rect 24977 -7267 25015 -7233
rect 25049 -7267 25087 -7233
rect 25121 -7267 25159 -7233
rect 25193 -7267 25231 -7233
rect 25265 -7267 25303 -7233
rect 25337 -7267 25375 -7233
rect 25409 -7267 25447 -7233
rect 25481 -7267 25519 -7233
rect 25553 -7267 25591 -7233
rect 25625 -7267 25663 -7233
rect 25697 -7267 25735 -7233
rect 25769 -7267 25807 -7233
rect 25841 -7267 25879 -7233
rect 25913 -7267 25951 -7233
rect 25985 -7267 26023 -7233
rect 26057 -7267 26095 -7233
rect 26129 -7267 26167 -7233
rect 26201 -7267 26239 -7233
rect 26273 -7267 26311 -7233
rect 26345 -7267 26383 -7233
rect 26417 -7267 26455 -7233
rect 26489 -7267 26527 -7233
rect 26561 -7267 26599 -7233
rect 26633 -7267 26671 -7233
rect 26705 -7267 26743 -7233
rect 26777 -7267 26815 -7233
rect 26849 -7267 26887 -7233
rect 26921 -7267 26959 -7233
rect 26993 -7267 27031 -7233
rect 27065 -7267 27103 -7233
rect 27137 -7267 27175 -7233
rect 27209 -7267 27247 -7233
rect 27281 -7267 27319 -7233
rect 27353 -7267 27391 -7233
rect 27425 -7267 27463 -7233
rect 27497 -7267 27535 -7233
rect 27569 -7267 27607 -7233
rect 27641 -7267 27679 -7233
rect 27713 -7267 27751 -7233
rect 27785 -7267 27823 -7233
rect 27857 -7267 27895 -7233
rect 27929 -7267 27967 -7233
rect 28001 -7267 28039 -7233
rect 28073 -7267 28111 -7233
rect 28145 -7267 28183 -7233
rect 28217 -7267 28255 -7233
rect 28289 -7267 28327 -7233
rect 28361 -7267 28399 -7233
rect 28433 -7267 28471 -7233
rect 28505 -7267 28543 -7233
rect 28577 -7267 28615 -7233
rect 28649 -7267 28687 -7233
rect 28721 -7267 28759 -7233
rect 28793 -7267 28831 -7233
rect 28865 -7267 28903 -7233
rect 28937 -7267 28975 -7233
rect 29009 -7267 29047 -7233
rect 29081 -7267 29119 -7233
rect 29153 -7267 29191 -7233
rect 29225 -7267 29263 -7233
rect 29297 -7267 29335 -7233
rect 29369 -7267 29407 -7233
rect 29441 -7267 29479 -7233
rect 29513 -7267 29551 -7233
rect 29585 -7267 29623 -7233
rect 29657 -7267 29695 -7233
rect 29729 -7267 29767 -7233
rect 29801 -7267 29839 -7233
rect 29873 -7267 29911 -7233
rect 29945 -7267 29983 -7233
rect 30017 -7267 30055 -7233
rect 30089 -7267 30127 -7233
rect 30161 -7267 30199 -7233
rect 30233 -7267 30271 -7233
rect 30305 -7267 30343 -7233
rect 30377 -7267 30415 -7233
rect 30449 -7267 30487 -7233
rect 30521 -7267 30559 -7233
rect 30593 -7267 30631 -7233
rect 30665 -7267 30703 -7233
rect 30737 -7267 30775 -7233
rect 30809 -7267 30847 -7233
rect 30881 -7267 30919 -7233
rect 30953 -7267 30991 -7233
rect 31025 -7267 31063 -7233
rect 31097 -7267 31135 -7233
rect 31169 -7267 31207 -7233
rect 31241 -7267 31279 -7233
rect 31313 -7267 31351 -7233
rect 31385 -7267 31423 -7233
rect 31457 -7267 31495 -7233
rect 31529 -7267 31567 -7233
rect 31601 -7267 31639 -7233
rect 31673 -7267 31711 -7233
rect 31745 -7267 31783 -7233
rect 31817 -7267 31855 -7233
rect 31889 -7267 31927 -7233
rect 31961 -7267 31999 -7233
rect 32033 -7267 32071 -7233
rect 32105 -7267 32143 -7233
rect 32177 -7267 32215 -7233
rect 32249 -7267 32287 -7233
rect 32321 -7267 32359 -7233
rect 32393 -7267 32431 -7233
rect 32465 -7267 32503 -7233
rect 32537 -7267 32575 -7233
rect 32609 -7267 32647 -7233
rect 32681 -7267 32719 -7233
rect 32753 -7267 32791 -7233
rect 32825 -7267 32863 -7233
rect 32897 -7267 32935 -7233
rect 32969 -7267 33007 -7233
rect 33041 -7267 33079 -7233
rect 33113 -7267 33151 -7233
rect 33185 -7267 33223 -7233
rect 33257 -7267 33295 -7233
rect 33329 -7267 33367 -7233
rect 33401 -7267 33439 -7233
rect 33473 -7267 33511 -7233
rect 33545 -7267 33583 -7233
rect 33617 -7267 33655 -7233
rect 33689 -7267 33727 -7233
rect 33761 -7267 33799 -7233
rect 33833 -7267 33871 -7233
rect 33905 -7267 33943 -7233
rect 33977 -7267 34015 -7233
rect 34049 -7267 34087 -7233
rect 34121 -7267 34159 -7233
rect 34193 -7267 34231 -7233
rect 34265 -7267 34303 -7233
rect 34337 -7267 34375 -7233
rect 34409 -7267 34447 -7233
rect 34481 -7267 34519 -7233
rect 34553 -7267 34591 -7233
rect 34625 -7267 34663 -7233
rect 34697 -7267 34735 -7233
rect 34769 -7267 34807 -7233
rect 34841 -7267 34879 -7233
rect 34913 -7267 34951 -7233
rect 34985 -7267 35023 -7233
rect 35057 -7267 35095 -7233
rect 35129 -7267 35167 -7233
rect 35201 -7267 35400 -7233
rect -17500 -7300 35400 -7267
<< metal2 >>
rect 300 360 17600 420
use XM_output_mirr_combined  XM_output_mirr_combined_0
timestamp 1663011646
transform 1 0 0 0 1 0
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_1
timestamp 1663011646
transform 1 0 0 0 1 7400
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_2
timestamp 1663011646
transform 1 0 0 0 1 -7400
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_3
timestamp 1663011646
transform 1 0 -17600 0 1 7400
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_4
timestamp 1663011646
transform 1 0 -17600 0 1 0
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_5
timestamp 1663011646
transform 1 0 -17600 0 1 -7400
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_6
timestamp 1663011646
transform 1 0 17600 0 1 7400
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_7
timestamp 1663011646
transform 1 0 17600 0 1 0
box 74 74 17826 7526
use XM_output_mirr_combined  XM_output_mirr_combined_8
timestamp 1663011646
transform 1 0 17600 0 1 -7400
box 74 74 17826 7526
<< end >>
