magic
tech sky130A
magscale 1 2
timestamp 1663029804
<< locali >>
rect 33895 33140 34005 33155
rect 33895 33085 33910 33140
rect 33990 33085 34005 33140
rect 33895 33070 34005 33085
rect 55194 32310 55348 32350
rect 33260 32140 33380 32155
rect 33260 32000 33275 32140
rect 33365 32000 33380 32140
rect 33260 31990 33380 32000
rect 52140 31560 52255 31580
rect 36440 31200 36900 31220
rect 36440 31140 36460 31200
rect 36880 31140 36900 31200
rect 52140 31190 52150 31560
rect 52240 31190 52255 31560
rect 52140 31175 52255 31190
rect 36440 31120 36900 31140
rect 55184 29702 55338 29742
rect 55174 27882 55328 27922
rect 52135 26440 52250 26455
rect 52135 26065 52145 26440
rect 52235 26065 52250 26440
rect 52135 26050 52250 26065
rect 34160 25810 36370 25850
rect 36420 25580 36940 25590
rect 33670 25570 36940 25580
rect 33670 25540 36430 25570
rect 36420 25530 36430 25540
rect 36930 25530 36940 25570
rect 36420 25510 36940 25530
rect 55178 25280 55332 25320
rect 32925 24465 33320 24480
rect 32925 24380 32940 24465
rect 33300 24380 33320 24465
rect 32925 24370 33320 24380
<< viali >>
rect 33910 33085 33990 33140
rect 33275 32000 33365 32140
rect 36460 31140 36880 31200
rect 52150 31190 52240 31560
rect 52145 26065 52235 26440
rect 36430 25530 36930 25570
rect 32940 24380 33300 24465
<< metal1 >>
rect 46750 37650 46800 38020
rect 46210 37580 46800 37650
rect 33895 33140 34005 33155
rect 33895 33085 33910 33140
rect 33990 33085 34005 33140
rect 33895 33070 34005 33085
rect 33475 32875 33520 33000
rect 33590 32990 33665 33000
rect 33590 32935 33600 32990
rect 33655 32935 33665 32990
rect 33590 32925 33665 32935
rect 33455 32865 33530 32875
rect 33455 32810 33465 32865
rect 33520 32810 33530 32865
rect 33455 32800 33530 32810
rect 33605 32800 33650 32925
rect 33730 32875 33775 33000
rect 33845 32990 33920 33000
rect 33845 32935 33855 32990
rect 33910 32935 33920 32990
rect 33845 32925 33920 32935
rect 33715 32865 33790 32875
rect 33715 32810 33725 32865
rect 33780 32810 33790 32865
rect 33715 32800 33790 32810
rect 33860 32800 33905 32925
rect 33520 32745 33865 32755
rect 33520 32715 33790 32745
rect 33780 32690 33790 32715
rect 33855 32690 33865 32745
rect 33780 32210 33865 32690
rect 36090 32690 36320 32760
rect 46210 32690 46280 37580
rect 47720 36710 47775 37940
rect 48190 36710 48240 38290
rect 47700 36700 47790 36710
rect 47700 36510 47710 36700
rect 47780 36510 47790 36700
rect 47700 36500 47790 36510
rect 48170 36700 48260 36710
rect 48170 36510 48180 36700
rect 48250 36510 48260 36700
rect 48170 36500 48260 36510
rect 33260 32140 33380 32155
rect 33260 32000 33275 32140
rect 33365 32000 33380 32140
rect 33260 31990 33380 32000
rect 35740 30980 35980 31000
rect 35740 30640 35760 30980
rect 35580 30630 35760 30640
rect 35960 30630 35980 30980
rect 35580 30580 35980 30630
rect 35761 27556 35862 27557
rect 35620 27495 35862 27556
rect 35761 27017 35862 27495
rect 35761 26613 35774 27017
rect 35848 26613 35862 27017
rect 35761 26603 35862 26613
rect 36090 25345 36160 32690
rect 36440 31200 36900 31220
rect 36440 31120 36460 31200
rect 36880 31120 36900 31200
rect 46335 31170 46440 31580
rect 36440 31100 36900 31120
rect 50680 31080 50730 37490
rect 57390 36205 57750 36265
rect 59485 36205 59860 36265
rect 61580 36205 61955 36265
rect 63670 36205 64910 36265
rect 57365 35845 57745 35905
rect 59490 35845 59865 35905
rect 61585 35845 61960 35905
rect 63690 35845 64655 35905
rect 57355 35305 57730 35365
rect 59465 35305 59840 35365
rect 61595 35305 61970 35365
rect 63660 35305 64405 35365
rect 57380 34715 57755 34775
rect 59460 34715 59835 34775
rect 61570 34715 61945 34775
rect 63655 34715 64140 34775
rect 57385 33805 57760 33865
rect 59460 33805 59835 33865
rect 61555 33805 61930 33865
rect 63700 33805 63905 33865
rect 52140 31560 52255 31580
rect 52140 31190 52150 31560
rect 52240 31190 52255 31560
rect 52140 31175 52255 31190
rect 55108 31074 56370 31134
rect 56292 31042 56370 31074
rect 56290 26556 56366 26586
rect 55094 26496 56366 26556
rect 52135 26440 52250 26455
rect 52135 26065 52145 26440
rect 52235 26065 52250 26440
rect 52135 26050 52250 26065
rect 36420 25570 36940 25590
rect 36420 25480 36430 25570
rect 36930 25480 36940 25570
rect 36420 25470 36940 25480
rect 36045 25335 36160 25345
rect 36045 25030 36055 25335
rect 36145 25030 36160 25335
rect 36045 25020 36160 25030
rect 32925 24465 33320 24480
rect 32925 24380 32940 24465
rect 33300 24380 33320 24465
rect 32925 24370 33320 24380
rect 36090 24050 36160 25020
rect 36090 23980 36400 24050
rect 63845 23825 63905 33805
rect 57370 23765 57745 23825
rect 59445 23765 59820 23825
rect 61580 23765 61955 23825
rect 63585 23765 63905 23825
rect 64080 22915 64140 34715
rect 57350 22855 57725 22915
rect 59460 22855 59835 22915
rect 61575 22855 61950 22915
rect 63635 22855 64140 22915
rect 64345 22325 64405 35305
rect 57370 22265 57745 22325
rect 59460 22265 59835 22325
rect 61575 22265 61950 22325
rect 63645 22265 64405 22325
rect 64595 21785 64655 35845
rect 57370 21725 57745 21785
rect 59475 21725 59850 21785
rect 61565 21725 61940 21785
rect 63700 21725 64655 21785
rect 64850 21425 64910 36205
rect 57360 21365 57735 21425
rect 59480 21365 59855 21425
rect 61570 21365 61945 21425
rect 63690 21365 64910 21425
<< via1 >>
rect 33910 33085 33990 33140
rect 33600 32935 33655 32990
rect 33465 32810 33520 32865
rect 33855 32935 33910 32990
rect 33725 32810 33780 32865
rect 33790 32690 33855 32745
rect 47710 36510 47780 36700
rect 48180 36510 48250 36700
rect 33275 32000 33365 32140
rect 35760 30630 35960 30980
rect 35774 26613 35848 27017
rect 36460 31140 36880 31180
rect 36460 31120 36880 31140
rect 52150 31190 52240 31560
rect 52145 26065 52235 26440
rect 36430 25530 36930 25540
rect 36430 25480 36930 25530
rect 36055 25030 36145 25335
rect 32940 24380 33300 24465
<< metal2 >>
rect 54790 37160 63285 37200
rect 54790 36800 54810 37160
rect 47700 36700 47790 36710
rect 47700 36510 47710 36700
rect 47780 36510 47790 36700
rect 47700 36500 47790 36510
rect 48170 36700 48260 36710
rect 48170 36510 48180 36700
rect 48250 36510 48260 36700
rect 54785 36620 54810 36800
rect 55190 36620 63285 37160
rect 54785 36600 63285 36620
rect 48170 36500 48260 36510
rect 55046 36460 55170 36462
rect 34240 36435 45110 36460
rect 34240 36045 34260 36435
rect 34515 36430 45110 36435
rect 34515 36060 45040 36430
rect 34515 36045 45110 36060
rect 34240 36020 45110 36045
rect 53625 35650 53690 36025
rect 56445 36130 56915 36600
rect 58545 36160 59040 36600
rect 58725 36145 58940 36160
rect 60650 36070 61180 36600
rect 62740 36095 63285 36600
rect 62640 36090 63285 36095
rect 54350 35650 54895 36025
rect 53625 35585 54895 35650
rect 33900 33140 34000 33145
rect 33900 33125 33910 33140
rect 33455 33085 33910 33125
rect 33990 33125 34000 33140
rect 33990 33110 34520 33125
rect 33990 33085 34210 33110
rect 33455 32990 34210 33085
rect 33455 32935 33600 32990
rect 33655 32935 33855 32990
rect 33910 32940 34210 32990
rect 34495 32940 34520 33110
rect 33910 32935 34520 32940
rect 33455 32925 34520 32935
rect 53710 33050 54520 35585
rect 33045 32865 33910 32875
rect 33045 32810 33465 32865
rect 33520 32810 33725 32865
rect 33780 32810 33910 32865
rect 33045 32745 33910 32810
rect 33045 32690 33790 32745
rect 33855 32690 33910 32745
rect 33045 32675 33910 32690
rect 53710 32715 55650 33050
rect 53710 32240 55996 32715
rect 55432 32200 55996 32240
rect 33260 32140 33380 32155
rect 33260 32000 33275 32140
rect 33365 32000 33380 32140
rect 33260 31990 33380 32000
rect 36440 31180 36900 31200
rect 36440 31120 36460 31180
rect 36880 31120 36900 31180
rect 36440 31100 36900 31120
rect 35740 30980 35980 31000
rect 35740 30630 35760 30980
rect 35960 30630 35980 30980
rect 35740 30610 35980 30630
rect 35760 27017 45180 27030
rect 35760 26613 35774 27017
rect 35848 26613 45180 27017
rect 35760 26600 45180 26613
rect 36420 25540 36940 25560
rect 36420 25480 36430 25540
rect 36930 25480 36940 25540
rect 36420 25470 36940 25480
rect 34665 25335 36160 25345
rect 34665 25030 36055 25335
rect 36145 25030 36160 25335
rect 34665 25020 36160 25030
rect 53900 24570 55890 25380
rect 53900 22045 54710 24570
rect 53600 21990 54895 22045
rect 53600 21605 53680 21990
rect 54610 21605 54895 21990
rect 56480 21035 56980 21530
rect 58550 21035 59100 21550
rect 60630 21035 61195 21540
rect 62895 21440 63110 21475
rect 62745 21035 63295 21440
rect 54785 21030 63295 21035
rect 54780 21020 63295 21030
rect 54780 20510 54810 21020
rect 55230 20510 63295 21020
rect 54780 20430 63295 20510
<< via2 >>
rect 43710 37930 44220 38270
rect 47710 36510 47780 36700
rect 48180 36510 48250 36700
rect 54810 36620 55190 37160
rect 34260 36045 34515 36435
rect 45040 36060 45430 36430
rect 53690 35650 54350 36390
rect 34210 32940 34495 33110
rect 54804 31204 55168 31558
rect 36460 31120 36880 31180
rect 35760 30630 35960 30980
rect 54882 26420 55210 26422
rect 54840 26090 55210 26420
rect 36430 25480 36930 25540
rect 53680 21230 54610 21990
rect 54810 20510 55230 21020
<< metal3 >>
rect 43670 38270 44270 38310
rect 43670 37930 43710 38270
rect 44220 37930 44270 38270
rect 34190 36435 34635 36460
rect 34190 36430 34260 36435
rect 34515 36430 34635 36435
rect 34190 36060 34230 36430
rect 34590 36060 34635 36430
rect 34190 36045 34260 36060
rect 34515 36045 34635 36060
rect 34190 36020 34635 36045
rect 34190 33110 34540 36020
rect 34190 32940 34210 33110
rect 34495 32940 34540 33110
rect 34190 32330 34540 32940
rect 34240 32200 34540 32330
rect 36410 32470 36940 32500
rect 43670 32470 44270 37930
rect 45000 36430 45470 38130
rect 54790 37160 55250 37200
rect 54790 36795 54810 37160
rect 47220 36700 47790 36710
rect 47220 36510 47710 36700
rect 47780 36510 47790 36700
rect 47220 36500 47790 36510
rect 48170 36700 49720 36710
rect 48170 36510 48180 36700
rect 48250 36510 49720 36700
rect 48170 36500 49720 36510
rect 54785 36620 54810 36795
rect 55190 36620 55250 37160
rect 45000 36060 45040 36430
rect 45430 36060 45470 36430
rect 45000 36020 45470 36060
rect 53612 36390 54420 36468
rect 53612 35650 53690 36390
rect 54350 35650 54420 36390
rect 53612 35578 54420 35650
rect 54785 36060 54840 36620
rect 55180 36060 55250 36620
rect 56840 37160 57650 37800
rect 56840 36660 56940 37160
rect 57560 36660 57650 37160
rect 56840 36590 57650 36660
rect 36410 32460 44270 32470
rect 36410 31920 36480 32460
rect 36880 31920 44270 32460
rect 36410 31880 44270 31920
rect 36410 31320 36940 31880
rect 54785 31578 55250 36060
rect 54785 31576 56340 31578
rect 54782 31558 56340 31576
rect 54782 31204 54804 31558
rect 55168 31204 56340 31558
rect 36440 31180 36900 31200
rect 36440 31120 36460 31180
rect 36880 31120 36900 31180
rect 54782 31176 56340 31204
rect 36440 31100 36900 31120
rect 35740 30980 35980 31000
rect 35740 30630 35760 30980
rect 35960 30630 35980 30980
rect 35740 30610 35980 30630
rect 57480 29855 57720 30020
rect 61085 30195 62590 30270
rect 59300 29670 59610 29800
rect 61085 29810 61855 30195
rect 62520 29810 62590 30195
rect 59755 29670 59780 29800
rect 61085 29785 62590 29810
rect 59300 29490 59780 29670
rect 56407 27820 56420 28090
rect 55650 27750 55670 27770
rect 61090 27800 62625 27835
rect 61090 27385 61850 27800
rect 62590 27385 62625 27800
rect 61090 27360 62625 27385
rect 54790 26456 55260 26460
rect 54790 26422 56470 26456
rect 54790 26420 54882 26422
rect 54790 26090 54840 26420
rect 55210 26090 56470 26422
rect 54790 26060 56470 26090
rect 54795 26054 56470 26060
rect 33845 24620 36555 24695
rect 33845 24140 34550 24620
rect 35760 24140 36555 24620
rect 33845 24090 36555 24140
rect 54795 23560 55260 26054
rect 54795 22580 54850 23560
rect 55150 22580 55260 23560
rect 53610 21990 54670 22040
rect 53610 21230 53680 21990
rect 54610 21230 54670 21990
rect 53610 21170 54670 21230
rect 54795 21020 55260 22580
rect 54795 20845 54810 21020
rect 54800 20510 54810 20845
rect 55230 20510 55260 21020
rect 54800 20430 55260 20510
<< via3 >>
rect 34230 36060 34260 36430
rect 34260 36060 34515 36430
rect 34515 36060 34590 36430
rect 54840 36620 55180 37130
rect 45040 36060 45430 36430
rect 53690 35650 54350 36390
rect 54840 36060 55180 36620
rect 56940 36660 57560 37160
rect 36480 31920 36880 32460
rect 35760 30630 35960 30980
rect 55465 29875 55925 30220
rect 57735 29855 58240 30245
rect 59610 29670 59755 30060
rect 61855 29810 62520 30195
rect 55465 27385 55950 27750
rect 57710 27380 58235 27765
rect 59620 27555 59860 28120
rect 61850 27385 62590 27800
rect 54840 26090 55200 26420
rect 34550 24140 35760 24620
rect 54850 22580 55150 23560
rect 53680 21230 54610 21990
<< metal4 >>
rect 52260 36470 52850 37560
rect 54780 37160 65400 37240
rect 54780 37130 56940 37160
rect 52260 36468 54190 36470
rect 34190 36430 34630 36460
rect 34190 36060 34230 36430
rect 34590 36060 34630 36430
rect 34190 36020 34630 36060
rect 45000 36430 45470 36460
rect 45000 36060 45040 36430
rect 45430 36060 45470 36430
rect 45000 36030 45470 36060
rect 52260 36390 54420 36468
rect 52260 35860 53690 36390
rect 53612 35650 53690 35860
rect 54350 35650 54420 36390
rect 54780 36060 54840 37130
rect 55180 36660 56940 37130
rect 57560 36660 65400 37160
rect 55180 36600 65400 36660
rect 55180 36060 55250 36600
rect 56840 36590 57650 36600
rect 54780 36000 55250 36060
rect 53612 35578 54420 35650
rect 36410 32460 36940 32500
rect 36410 31920 36480 32460
rect 36880 31920 36940 32460
rect 36410 31840 36940 31920
rect 35740 30980 36320 31000
rect 35740 30630 35760 30980
rect 35960 30630 36320 30980
rect 35740 30610 36320 30630
rect 61810 30435 62585 30475
rect 55435 30230 56170 30260
rect 55435 30220 55710 30230
rect 55435 29875 55465 30220
rect 56135 29920 56170 30230
rect 55925 29875 56170 29920
rect 55435 29850 56170 29875
rect 57695 30245 58260 30270
rect 57695 29855 57735 30245
rect 58240 29855 58260 30245
rect 61810 30195 62015 30435
rect 59865 30160 60165 30190
rect 59865 30095 59900 30160
rect 57695 29835 58260 29855
rect 59600 30060 59900 30095
rect 59600 29670 59610 30060
rect 59755 29920 59900 30060
rect 60140 29920 60165 30160
rect 59755 29895 60165 29920
rect 59755 29670 59775 29895
rect 61810 29810 61855 30195
rect 62555 29930 62585 30435
rect 62520 29810 62585 29930
rect 61810 29780 62585 29810
rect 59600 29655 59775 29670
rect 59600 28120 59885 28140
rect 55440 27750 56175 27820
rect 55440 27385 55465 27750
rect 55950 27705 56175 27750
rect 56125 27390 56175 27705
rect 55950 27385 56175 27390
rect 55440 27355 56175 27385
rect 57695 27765 58255 27790
rect 57695 27380 57710 27765
rect 58235 27380 58255 27765
rect 59600 27555 59620 28120
rect 59860 27735 59885 28120
rect 61810 27800 62620 27830
rect 59860 27715 60200 27735
rect 59860 27555 59905 27715
rect 59600 27510 59905 27555
rect 59885 27475 59905 27510
rect 60180 27475 60200 27715
rect 59885 27465 60200 27475
rect 57695 27360 58255 27380
rect 61810 27385 61850 27800
rect 62590 27385 62620 27800
rect 61810 27260 62015 27385
rect 62580 27260 62620 27385
rect 61810 27225 62620 27260
rect 54790 26420 55250 26460
rect 54790 26090 54840 26420
rect 55200 26090 55250 26420
rect 54790 26060 55250 26090
rect 34440 24620 35960 24700
rect 34440 24140 34550 24620
rect 35760 24140 35960 24620
rect 34440 23320 35960 24140
rect 54760 23560 55240 23630
rect 54760 22580 54850 23560
rect 55150 22580 55240 23560
rect 54760 22520 55240 22580
rect 53610 21990 54670 22040
rect 53610 21230 53680 21990
rect 54610 21230 54670 21990
rect 53610 21170 54670 21230
<< via4 >>
rect 34230 36060 34590 36430
rect 45040 36060 45430 36430
rect 53690 35650 54350 36390
rect 54840 36060 55180 37130
rect 56940 36660 57560 37160
rect 36480 31920 36880 32460
rect 55710 30220 56135 30230
rect 55710 29920 55925 30220
rect 55925 29920 56135 30220
rect 57735 29865 58240 30245
rect 62015 30195 62555 30435
rect 59900 29920 60140 30160
rect 62015 29930 62520 30195
rect 62520 29930 62555 30195
rect 55710 27390 55950 27705
rect 55950 27390 56125 27705
rect 57715 27385 58235 27765
rect 59905 27475 60180 27715
rect 62015 27385 62580 27700
rect 62015 27260 62580 27385
rect 54840 26090 55200 26420
rect 34550 24140 35760 24620
rect 54850 22580 55150 23560
rect 53680 21230 54610 21990
<< metal5 >>
rect 54780 37160 57650 37240
rect 54780 37130 56940 37160
rect 53612 36460 54420 36468
rect 34170 36430 54420 36460
rect 34170 36060 34230 36430
rect 34590 36060 45040 36430
rect 45430 36390 54420 36430
rect 45430 36060 53690 36390
rect 34170 35650 53690 36060
rect 54350 35650 54420 36390
rect 34170 35640 54420 35650
rect 53612 35578 54420 35640
rect 54780 36060 54840 37130
rect 55180 36660 56940 37130
rect 57560 36660 57650 37160
rect 55180 36590 57650 36660
rect 55180 36060 55330 36590
rect 36330 32460 37030 32510
rect 36330 31920 36480 32460
rect 36880 31920 37030 32460
rect 36330 24710 37030 31920
rect 34480 24620 37040 24710
rect 34480 24140 34550 24620
rect 35760 24140 37040 24620
rect 34480 24080 37040 24140
rect 53630 22040 54080 35578
rect 54780 35180 55330 36060
rect 54550 34620 55330 35180
rect 54550 26420 55250 34620
rect 57695 30245 58260 30270
rect 55705 29920 55710 30230
rect 57695 29865 57735 30245
rect 58240 29910 58260 30245
rect 59865 30190 59895 30215
rect 59865 30160 60165 30190
rect 59865 29920 59900 30160
rect 60140 29920 60165 30160
rect 58240 29865 58265 29910
rect 59865 29895 60165 29920
rect 57695 29835 58265 29865
rect 57685 27765 58260 27790
rect 57685 27385 57715 27765
rect 58235 27385 58260 27765
rect 59875 27715 60200 27740
rect 59875 27475 59905 27715
rect 60180 27475 60200 27715
rect 59875 27400 60200 27475
rect 57685 27360 58260 27385
rect 54550 26090 54840 26420
rect 55200 26090 55250 26420
rect 54550 23560 55250 26090
rect 54550 22580 54850 23560
rect 55150 22580 55250 23560
rect 54550 22520 55250 22580
rect 53610 21990 54670 22040
rect 53610 21230 53680 21990
rect 54610 21230 54670 21990
rect 53610 21170 54670 21230
use core_osc  X1
timestamp 1662665761
transform 1 0 46065 0 1 21045
box 9175 3425 16085 12111
use buffer_amp_vop  X3
timestamp 1662952744
transform 1 0 26070 0 1 10600
box 10225 10400 29180 26030
use cap_bank  X4
timestamp 1663029804
transform 1 0 52305 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X5
timestamp 1663029804
transform 1 0 54405 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X6
timestamp 1663029804
transform 1 0 52305 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X7
timestamp 1663029804
transform 1 0 54405 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X8
timestamp 1663029804
transform 1 0 56505 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X9
timestamp 1663029804
transform 1 0 58605 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X10
timestamp 1663029804
transform 1 0 56505 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X11
timestamp 1663029804
transform 1 0 58605 0 -1 34725
box 3300 -1540 5112 5514
use bias_calc  bias_calc_0
timestamp 1662665484
transform 1 0 14295 0 1 25060
box 16846 -965 21340 7275
use output_buffer  output_buffer_0
timestamp 1662517639
transform 1 0 34825 0 1 39195
box 8845 -1865 22825 2478
use sky130_fd_pr__pfet_01v8_lvt_75KH85  sky130_fd_pr__pfet_01v8_lvt_75KH85_0
timestamp 1662690363
transform 1 0 33689 0 1 32864
box -359 -284 359 284
<< labels >>
rlabel metal5 53630 21190 54080 36450 1 VDD
rlabel metal5 36330 24100 37030 32510 1 GND
rlabel metal1 64850 21365 64910 36265 1 CTRL1
rlabel metal1 64595 21725 64655 35905 1 CTRL2
rlabel metal1 64345 22265 64405 35365 1 CTRL3
rlabel metal1 64080 22855 64140 34775 1 CTRL4
rlabel metal1 63845 23765 63905 33865 1 CTRL5
rlabel metal2 60650 36070 61180 37200 1 GND
<< end >>
