magic
tech sky130A
magscale 1 2
timestamp 1662863789
<< locali >>
rect 24600 25950 24740 25990
rect 19760 21370 20200 21410
rect 24590 18790 24730 18830
rect 24590 17610 24730 17650
rect 19700 16820 20200 16860
rect 19750 15740 20210 15780
rect 19750 14940 20210 14980
rect 24590 10440 24730 10480
<< metal1 >>
rect 10240 22090 20210 22160
rect 20140 20480 20210 22090
rect 19740 19800 20080 19870
rect 20010 19200 20080 19800
rect 19990 19180 20100 19200
rect 19990 19100 20010 19180
rect 20080 19100 20100 19180
rect 19990 19080 20100 19100
rect 19700 19000 19910 19070
rect 19840 18650 19910 19000
rect 21660 18650 21770 18670
rect 19840 18580 21680 18650
rect 21750 18580 21770 18650
rect 21660 18560 21770 18580
rect 22120 18440 22230 18790
rect 22120 18380 22140 18440
rect 22210 18380 22230 18440
rect 22120 18360 22230 18380
rect 22820 18310 22930 18790
rect 26390 18750 26750 18800
rect 26650 18700 26750 18750
rect 26650 18640 26670 18700
rect 26730 18640 26750 18700
rect 26650 18620 26750 18640
rect 27350 18570 27450 18820
rect 27350 18510 27370 18570
rect 27430 18510 27450 18570
rect 27350 18490 27450 18510
rect 19750 17900 19820 18270
rect 22820 18250 22840 18310
rect 22910 18250 22930 18310
rect 22820 18230 22930 18250
rect 22120 18190 22230 18200
rect 22120 18110 22130 18190
rect 22220 18110 22230 18190
rect 21660 17900 21770 17920
rect 19750 17830 21680 17900
rect 21750 17830 21770 17900
rect 21660 17810 21770 17830
rect 22120 17610 22230 18110
rect 22820 18060 22930 18070
rect 22820 17980 22830 18060
rect 22920 17980 22930 18060
rect 22820 17610 22930 17980
rect 27350 17930 27450 17940
rect 27350 17850 27360 17930
rect 27440 17850 27450 17930
rect 26650 17800 26750 17810
rect 26650 17720 26660 17800
rect 26740 17720 26750 17800
rect 26650 17610 26750 17720
rect 27350 17610 27450 17850
rect 20130 17470 20240 17490
rect 19680 17400 20150 17470
rect 20220 17400 20240 17470
rect 20130 17380 20240 17400
rect 20140 13450 20202 15956
rect 10230 13380 20202 13450
<< via1 >>
rect 20010 19100 20080 19180
rect 21680 18580 21750 18650
rect 22140 18380 22210 18440
rect 26670 18640 26730 18700
rect 27370 18510 27430 18570
rect 22840 18250 22910 18310
rect 22130 18110 22220 18190
rect 21680 17830 21750 17900
rect 22830 17980 22920 18060
rect 27360 17850 27440 17930
rect 26660 17720 26740 17800
rect 20150 17400 20220 17470
<< metal2 >>
rect 18710 25420 20300 25860
rect 18710 20900 19000 25420
rect 19990 19180 20100 19200
rect 19990 19100 20010 19180
rect 20080 19100 20100 19180
rect 19990 19080 20100 19100
rect 22120 18700 29180 18720
rect 21660 18650 21770 18670
rect 21660 18580 21680 18650
rect 21750 18580 21770 18650
rect 22120 18640 26670 18700
rect 26730 18640 29180 18700
rect 22120 18620 29180 18640
rect 21660 18560 21770 18580
rect 22120 18570 29180 18590
rect 22120 18510 27370 18570
rect 27430 18510 29180 18570
rect 22120 18490 29180 18510
rect 22120 18440 29180 18460
rect 22120 18380 22140 18440
rect 22210 18380 29180 18440
rect 22120 18360 29180 18380
rect 22120 18310 29180 18330
rect 22120 18250 22840 18310
rect 22910 18250 29180 18310
rect 22120 18230 29180 18250
rect 22120 18190 29180 18200
rect 22120 18110 22130 18190
rect 22220 18110 29180 18190
rect 22120 18100 29180 18110
rect 22120 18060 29180 18070
rect 22120 17980 22830 18060
rect 22920 17980 29180 18060
rect 22120 17970 29180 17980
rect 22120 17930 29180 17940
rect 21660 17900 21770 17920
rect 21660 17830 21680 17900
rect 21750 17830 21770 17900
rect 22120 17850 27360 17930
rect 27440 17850 29180 17930
rect 22120 17840 29180 17850
rect 21660 17810 21770 17830
rect 22120 17800 29180 17810
rect 22120 17720 26660 17800
rect 26740 17720 29180 17800
rect 22120 17710 29180 17720
rect 20130 17470 20240 17490
rect 20130 17400 20150 17470
rect 20220 17400 20240 17470
rect 20130 17380 20240 17400
rect 17580 16990 19440 17020
rect 17580 16760 17610 16990
rect 17790 16760 19440 16990
rect 17580 16730 19440 16760
rect 10240 16000 19660 16430
rect 19230 15680 19660 16000
rect 17580 14390 18350 14420
rect 17580 14150 17610 14390
rect 17810 14150 18350 14390
rect 17580 14130 18350 14150
rect 19520 11010 19820 14420
rect 20650 13760 21050 15850
rect 20640 13470 21050 13760
rect 20640 13200 21040 13470
rect 20640 12840 20660 13200
rect 21010 12840 21040 13200
rect 20640 12820 21040 12840
rect 19520 10570 20250 11010
<< via2 >>
rect 20210 20620 20440 20930
rect 20010 19100 20080 19180
rect 21680 18580 21750 18650
rect 21680 17830 21750 17900
rect 20150 17400 20220 17470
rect 17610 16760 17790 16990
rect 17610 14150 17810 14390
rect 20660 12840 21010 13200
<< metal3 >>
rect 15670 20930 20500 20980
rect 15670 20620 20210 20930
rect 20440 20620 20500 20930
rect 15670 20580 20500 20620
rect 15670 20480 16440 20580
rect 15670 20270 16330 20480
rect 19990 19180 20410 19200
rect 19990 19100 20010 19180
rect 20080 19100 20410 19180
rect 19990 19080 20410 19100
rect 21150 18760 21450 26030
rect 22650 18670 22760 18830
rect 23350 18760 23650 26030
rect 21660 18650 22760 18670
rect 21660 18580 21680 18650
rect 21750 18580 22760 18650
rect 21660 18560 22760 18580
rect 25635 18330 25835 18939
rect 27680 18330 27880 18934
rect 19870 18100 27880 18330
rect 17540 16990 17840 17020
rect 17540 16760 17610 16990
rect 17790 16760 17840 16990
rect 10348 15604 10872 16712
rect 17540 14390 17840 16760
rect 17540 14150 17610 14390
rect 17810 14150 17840 14390
rect 17540 14130 17840 14150
rect 19870 13970 20070 18100
rect 21660 17900 22760 17920
rect 21660 17830 21680 17900
rect 21750 17830 22760 17900
rect 21660 17810 22760 17830
rect 20130 17470 20400 17490
rect 20130 17400 20150 17470
rect 20220 17400 20400 17470
rect 20130 17380 20400 17400
rect 19820 13570 20070 13970
rect 15850 13200 21040 13220
rect 15850 12840 20660 13200
rect 21010 12840 21040 13200
rect 15850 12820 21040 12840
rect 21150 10400 21450 17670
rect 22650 17570 22760 17810
rect 23350 10410 23650 17680
rect 25635 17490 25835 18100
rect 27680 17630 27880 18100
<< metal4 >>
rect 10225 20205 10250 20270
use buffer_amp  X1
timestamp 1662405622
transform 1 0 15140 0 1 17350
box 5000 1400 9520 8676
use buffer_amp  X2
timestamp 1662405622
transform 1 0 19660 0 -1 19081
box 5000 1400 9520 8676
use buffer_amp  X3
timestamp 1662405622
transform 1 0 15140 0 -1 19081
box 5000 1400 9520 8676
use buffer_amp  X4
timestamp 1662405622
transform 1 0 19660 0 1 17350
box 5000 1400 9520 8676
use amp_dec  X5
timestamp 1662519997
transform 0 1 9640 -1 0 26439
box 5000 590 10199 10196
use vop_dec  X6
timestamp 1662515827
transform 0 1 9830 -1 0 21409
box 5600 400 10899 9996
<< labels >>
rlabel metal2 10240 16000 19660 16430 1 VOP
rlabel metal3 15850 12820 20660 13220 1 GND
rlabel metal1 10230 13380 20140 13450 1 BIAS
rlabel metal3 21150 18760 21450 26030 1 OUT180
rlabel metal3 23350 18760 23650 26030 1 OUT0
rlabel metal3 21150 10400 21450 17670 1 OUT270
rlabel metal3 23350 10410 23650 17680 1 OUT90
rlabel locali 19760 21370 20200 21410 1 SUB
rlabel metal1 10240 22090 20210 22160 1 BIAS
rlabel space 10230 20009 11310 20399 1 AMP
rlabel metal4 10225 20205 10250 20270 1 AMP
rlabel metal2 26730 18620 29180 18720 1 I4B
rlabel metal2 27430 18490 29180 18590 1 I4A
rlabel metal2 22210 18360 29180 18460 1 I1B
rlabel metal2 22910 18230 29180 18330 1 I1A
rlabel metal2 26740 18100 29180 18200 1 I3B
rlabel metal2 27440 17970 29180 18070 1 I3A
rlabel metal2 22920 17840 29180 17940 1 I2A
rlabel metal2 22220 17710 29180 17810 1 I2B
rlabel metal2 19520 10570 19820 14420 1 VDD
<< end >>
