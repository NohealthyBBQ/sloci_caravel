magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -236 -319 236 319
<< nmos >>
rect -50 -181 50 119
<< ndiff >>
rect -108 88 -50 119
rect -108 54 -96 88
rect -62 54 -50 88
rect -108 20 -50 54
rect -108 -14 -96 20
rect -62 -14 -50 20
rect -108 -48 -50 -14
rect -108 -82 -96 -48
rect -62 -82 -50 -48
rect -108 -116 -50 -82
rect -108 -150 -96 -116
rect -62 -150 -50 -116
rect -108 -181 -50 -150
rect 50 88 108 119
rect 50 54 62 88
rect 96 54 108 88
rect 50 20 108 54
rect 50 -14 62 20
rect 96 -14 108 20
rect 50 -48 108 -14
rect 50 -82 62 -48
rect 96 -82 108 -48
rect 50 -116 108 -82
rect 50 -150 62 -116
rect 96 -150 108 -116
rect 50 -181 108 -150
<< ndiffc >>
rect -96 54 -62 88
rect -96 -14 -62 20
rect -96 -82 -62 -48
rect -96 -150 -62 -116
rect 62 54 96 88
rect 62 -14 96 20
rect 62 -82 96 -48
rect 62 -150 96 -116
<< psubdiff >>
rect -210 259 -85 293
rect -51 259 -17 293
rect 17 259 51 293
rect 85 259 210 293
rect -210 -259 -176 259
rect 176 -259 210 259
rect -210 -293 -85 -259
rect -51 -293 -17 -259
rect 17 -293 51 -259
rect 85 -293 210 -259
<< psubdiffcont >>
rect -85 259 -51 293
rect -17 259 17 293
rect 51 259 85 293
rect -85 -293 -51 -259
rect -17 -293 17 -259
rect 51 -293 85 -259
<< poly >>
rect -50 191 50 207
rect -50 157 -17 191
rect 17 157 50 191
rect -50 119 50 157
rect -50 -207 50 -181
<< polycont >>
rect -17 157 17 191
<< locali >>
rect -210 259 -85 293
rect -51 259 -17 293
rect 17 259 51 293
rect 85 259 210 293
rect -210 -259 -176 259
rect -50 157 -17 191
rect 17 157 50 191
rect -96 94 -62 123
rect -96 22 -62 54
rect -96 -48 -62 -14
rect -96 -116 -62 -84
rect -96 -185 -62 -156
rect 62 94 96 123
rect 62 22 96 54
rect 62 -48 96 -14
rect 62 -116 96 -84
rect 62 -185 96 -156
rect 176 -259 210 259
rect -210 -293 -85 -259
rect -51 -293 -17 -259
rect 17 -293 51 -259
rect 85 -293 210 -259
<< viali >>
rect -17 157 17 191
rect -96 88 -62 94
rect -96 60 -62 88
rect -96 20 -62 22
rect -96 -12 -62 20
rect -96 -82 -62 -50
rect -96 -84 -62 -82
rect -96 -150 -62 -122
rect -96 -156 -62 -150
rect 62 88 96 94
rect 62 60 96 88
rect 62 20 96 22
rect 62 -12 96 20
rect 62 -82 96 -50
rect 62 -84 96 -82
rect 62 -150 96 -122
rect 62 -156 96 -150
<< metal1 >>
rect -46 191 46 197
rect -46 157 -17 191
rect 17 157 46 191
rect -46 151 46 157
rect -102 94 -56 119
rect -102 60 -96 94
rect -62 60 -56 94
rect -102 22 -56 60
rect -102 -12 -96 22
rect -62 -12 -56 22
rect -102 -50 -56 -12
rect -102 -84 -96 -50
rect -62 -84 -56 -50
rect -102 -122 -56 -84
rect -102 -156 -96 -122
rect -62 -156 -56 -122
rect -102 -181 -56 -156
rect 56 94 102 119
rect 56 60 62 94
rect 96 60 102 94
rect 56 22 102 60
rect 56 -12 62 22
rect 96 -12 102 22
rect 56 -50 102 -12
rect 56 -84 62 -50
rect 96 -84 102 -50
rect 56 -122 102 -84
rect 56 -156 62 -122
rect 96 -156 102 -122
rect 56 -181 102 -156
<< properties >>
string FIXED_BBOX -193 -276 193 276
<< end >>
