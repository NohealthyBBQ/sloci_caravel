magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -349 -300 349 300
<< nmoslvt >>
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
<< ndiff >>
rect -221 85 -159 100
rect -221 51 -209 85
rect -175 51 -159 85
rect -221 17 -159 51
rect -221 -17 -209 17
rect -175 -17 -159 17
rect -221 -51 -159 -17
rect -221 -85 -209 -51
rect -175 -85 -159 -51
rect -221 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 221 100
rect 159 51 175 85
rect 209 51 221 85
rect 159 17 221 51
rect 159 -17 175 17
rect 209 -17 221 17
rect 159 -51 221 -17
rect 159 -85 175 -51
rect 209 -85 221 -51
rect 159 -100 221 -85
<< ndiffc >>
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
<< psubdiff >>
rect -323 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 323 274
rect -323 153 -289 240
rect -323 85 -289 119
rect 289 153 323 240
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect -323 -240 -289 -153
rect 289 -119 323 -85
rect 289 -240 323 -153
rect -323 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 323 -240
<< psubdiffcont >>
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect -323 119 -289 153
rect 289 119 323 153
rect -323 51 -289 85
rect -323 -17 -289 17
rect -323 -85 -289 -51
rect 289 51 323 85
rect 289 -17 323 17
rect 289 -85 323 -51
rect -323 -153 -289 -119
rect 289 -153 323 -119
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
<< poly >>
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 129 100 159 122
rect -159 -122 -129 -100
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
<< polycont >>
rect -65 138 -31 172
rect 127 138 161 172
rect -161 -172 -127 -138
rect 31 -172 65 -138
<< locali >>
rect -323 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 323 274
rect -323 153 -289 240
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 289 153 323 240
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect -323 -119 -289 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect 289 -119 323 -85
rect -323 -240 -289 -153
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 289 -240 323 -153
rect -323 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 323 -240
<< viali >>
rect -65 138 -31 172
rect 127 138 161 172
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect -161 -172 -127 -138
rect 31 -172 65 -138
<< metal1 >>
rect -77 175 -19 178
rect 115 175 173 178
rect -90 172 175 175
rect -90 140 -65 172
rect -77 138 -65 140
rect -31 140 127 172
rect -31 138 -19 140
rect -77 132 -19 138
rect 115 138 127 140
rect 161 140 175 172
rect 161 138 173 140
rect 115 132 173 138
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect -173 -138 -115 -132
rect -173 -140 -161 -138
rect -175 -172 -161 -140
rect -127 -140 -115 -138
rect 19 -138 77 -132
rect 19 -140 31 -138
rect -127 -172 31 -140
rect 65 -140 77 -138
rect 65 -172 80 -140
rect -175 -175 80 -172
rect -173 -178 -115 -175
rect 19 -178 77 -175
<< properties >>
string FIXED_BBOX -306 -257 306 257
<< end >>
