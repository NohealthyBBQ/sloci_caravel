magic
tech sky130A
timestamp 1663011646
<< locali >>
rect 300 1600 3000 1650
rect 300 950 1410 1000
rect 1840 950 3000 1000
rect 300 300 3000 350
<< metal1 >>
rect 1545 1036 1705 1050
rect 1545 914 1564 1036
rect 1686 914 1705 1036
rect 1545 900 1705 914
<< via1 >>
rect 1564 914 1686 1036
<< metal2 >>
rect 1550 1036 1700 1055
rect 1550 914 1564 1036
rect 1686 914 1700 1036
rect 1550 895 1700 914
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0
array 0 4 644 0 2 644
timestamp 1663011646
transform 1 0 0 0 1 0
box 0 0 670 670
<< end >>
