magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -8726 10225 -8100 11452
<< locali >>
rect -10880 11217 -10820 11240
rect -10880 11183 -10867 11217
rect -10833 11183 -10820 11217
rect -10880 11145 -10820 11183
rect -10880 11111 -10867 11145
rect -10833 11111 -10820 11145
rect -10880 11073 -10820 11111
rect -10880 11039 -10867 11073
rect -10833 11039 -10820 11073
rect -10880 11001 -10820 11039
rect -10880 10967 -10867 11001
rect -10833 10967 -10820 11001
rect -10880 10929 -10820 10967
rect -10880 10895 -10867 10929
rect -10833 10895 -10820 10929
rect -10880 10857 -10820 10895
rect -10880 10823 -10867 10857
rect -10833 10823 -10820 10857
rect -10880 10785 -10820 10823
rect -10880 10751 -10867 10785
rect -10833 10751 -10820 10785
rect -10880 10713 -10820 10751
rect -10880 10679 -10867 10713
rect -10833 10679 -10820 10713
rect -10880 10641 -10820 10679
rect -10880 10607 -10867 10641
rect -10833 10607 -10820 10641
rect -10880 10569 -10820 10607
rect -10880 10535 -10867 10569
rect -10833 10535 -10820 10569
rect -10880 10497 -10820 10535
rect -10880 10463 -10867 10497
rect -10833 10463 -10820 10497
rect -10880 10425 -10820 10463
rect -10880 10391 -10867 10425
rect -10833 10391 -10820 10425
rect -10880 10353 -10820 10391
rect -10880 10319 -10867 10353
rect -10833 10319 -10820 10353
rect -10880 10281 -10820 10319
rect -10880 10247 -10867 10281
rect -10833 10247 -10820 10281
rect -10880 10209 -10820 10247
rect -10880 10175 -10867 10209
rect -10833 10175 -10820 10209
rect -8800 10551 -8680 10580
rect -8800 10229 -8793 10551
rect -8687 10229 -8680 10551
rect -8800 10200 -8680 10229
rect -10880 10137 -10820 10175
rect -10880 10103 -10867 10137
rect -10833 10103 -10820 10137
rect -10880 10080 -10820 10103
rect -6920 9900 -6780 10760
rect -1960 10660 4480 10940
rect -1960 10600 1560 10660
rect -2980 9253 -2820 9280
rect -2980 9147 -2953 9253
rect -2847 9147 -2820 9253
rect -2980 8990 -2820 9147
rect -3350 8950 -1990 8990
rect -7740 8580 -7620 8860
rect -3330 8480 -2030 8490
rect -3350 8450 -1960 8480
rect -9000 8140 -8880 8440
rect -14000 7490 -13900 8080
rect -10900 7490 -10800 8080
rect -14030 7480 -10800 7490
rect -2040 6400 -1940 6840
rect -860 6400 -660 6820
rect 440 6400 640 6820
rect 1720 6400 1920 6820
rect 3020 6400 3220 6820
rect 4300 6400 4400 6860
rect 4620 333 5080 400
rect 4620 227 4689 333
rect 5011 227 5080 333
rect 4620 180 5080 227
rect 4560 -40 9140 20
rect 4560 -220 9140 -160
rect 4560 -580 9140 -520
rect 4580 -960 6100 -900
rect 7600 -960 9120 -900
rect 4560 -1140 6100 -1080
rect 7620 -1140 9140 -1080
rect 4580 -1500 6100 -1440
rect 7620 -1480 9140 -1420
rect 4560 -1880 9140 -1820
rect 4560 -2060 9140 -2000
rect -2120 -2400 -1960 -2380
rect -2120 -2427 4360 -2400
rect 4560 -2420 9140 -2360
rect -2120 -2533 -1553 -2427
rect -1447 -2480 4360 -2427
rect -1447 -2533 4400 -2480
rect -2120 -2580 4400 -2533
rect -2120 -2600 -1860 -2580
rect 4300 -2780 4400 -2580
rect 8480 -2780 9420 -2740
rect 9620 -2847 9920 -2840
rect 9620 -2953 9645 -2847
rect 9895 -2953 9920 -2847
rect 9620 -2960 9920 -2953
rect 33500 -2847 33800 -2840
rect 33500 -2953 33525 -2847
rect 33775 -2953 33800 -2847
rect 33500 -2960 33800 -2953
rect 61800 -2847 62100 -2840
rect 61800 -2953 61825 -2847
rect 62075 -2953 62100 -2847
rect 61800 -2960 62100 -2953
rect 7700 -3420 9500 -3260
rect -14180 -3820 -13640 -3520
rect 7700 -3960 9500 -3840
rect -14200 -10160 -13640 -9020
rect 8100 -10296 9500 -10200
<< viali >>
rect -10867 11183 -10833 11217
rect -10867 11111 -10833 11145
rect -10867 11039 -10833 11073
rect -10867 10967 -10833 11001
rect -10867 10895 -10833 10929
rect -10867 10823 -10833 10857
rect -10867 10751 -10833 10785
rect -10867 10679 -10833 10713
rect -10867 10607 -10833 10641
rect -10867 10535 -10833 10569
rect -10867 10463 -10833 10497
rect -10867 10391 -10833 10425
rect -10867 10319 -10833 10353
rect -10867 10247 -10833 10281
rect -10867 10175 -10833 10209
rect -8793 10229 -8687 10551
rect -10867 10103 -10833 10137
rect -2953 9147 -2847 9253
rect 4689 227 5011 333
rect -1553 -2533 -1447 -2427
rect 9645 -2953 9895 -2847
rect 33525 -2953 33775 -2847
rect 61825 -2953 62075 -2847
<< metal1 >>
rect -10910 11230 -10790 11260
rect -10910 11178 -10876 11230
rect -10824 11178 -10790 11230
rect -10910 11166 -10790 11178
rect -10910 11114 -10876 11166
rect -10824 11114 -10790 11166
rect 1190 11176 1310 11200
rect 1190 11124 1224 11176
rect 1276 11124 1310 11176
rect -10910 11111 -10867 11114
rect -10833 11111 -10790 11114
rect -10910 11102 -10790 11111
rect -10910 11050 -10876 11102
rect -10824 11050 -10790 11102
rect -10910 11039 -10867 11050
rect -10833 11039 -10790 11050
rect -7750 11106 -7670 11120
rect -7750 11054 -7736 11106
rect -7684 11054 -7670 11106
rect 1190 11100 1310 11124
rect -7750 11040 -7670 11054
rect -10910 11038 -10790 11039
rect -10910 10986 -10876 11038
rect -10824 10986 -10790 11038
rect -10910 10974 -10867 10986
rect -10833 10974 -10790 10986
rect -10910 10922 -10876 10974
rect -10824 10922 -10790 10974
rect -10910 10910 -10867 10922
rect -10833 10910 -10790 10922
rect -10910 10858 -10876 10910
rect -10824 10858 -10790 10910
rect -10910 10857 -10790 10858
rect -10910 10846 -10867 10857
rect -10833 10846 -10790 10857
rect -10910 10794 -10876 10846
rect -10824 10794 -10790 10846
rect -10910 10785 -10790 10794
rect -10910 10782 -10867 10785
rect -10833 10782 -10790 10785
rect -10910 10730 -10876 10782
rect -10824 10730 -10790 10782
rect -10910 10718 -10790 10730
rect -10910 10666 -10876 10718
rect -10824 10666 -10790 10718
rect -10910 10654 -10790 10666
rect -10910 10602 -10876 10654
rect -10824 10602 -10790 10654
rect -10910 10590 -10790 10602
rect -10910 10538 -10876 10590
rect -10824 10538 -10790 10590
rect -10910 10535 -10867 10538
rect -10833 10535 -10790 10538
rect -10910 10526 -10790 10535
rect -10910 10474 -10876 10526
rect -10824 10474 -10790 10526
rect -10910 10463 -10867 10474
rect -10833 10463 -10790 10474
rect -10910 10462 -10790 10463
rect -10910 10410 -10876 10462
rect -10824 10410 -10790 10462
rect -10910 10398 -10867 10410
rect -10833 10398 -10790 10410
rect -10910 10346 -10876 10398
rect -10824 10346 -10790 10398
rect -10910 10334 -10867 10346
rect -10833 10334 -10790 10346
rect -10910 10282 -10876 10334
rect -10824 10282 -10790 10334
rect -10910 10281 -10790 10282
rect -10910 10270 -10867 10281
rect -10833 10270 -10790 10281
rect -10910 10218 -10876 10270
rect -10824 10218 -10790 10270
rect -10910 10209 -10790 10218
rect -10910 10206 -10867 10209
rect -10833 10206 -10790 10209
rect -10910 10154 -10876 10206
rect -10824 10154 -10790 10206
rect -10910 10142 -10790 10154
rect -10910 10090 -10876 10142
rect -10824 10090 -10790 10142
rect -10910 10060 -10790 10090
rect -11458 9858 -10653 9906
rect -10600 8810 -10540 11000
rect -8806 10580 -8674 10592
rect -8810 10576 -8670 10580
rect -8810 10204 -8798 10576
rect -8682 10204 -8670 10576
rect -8230 10566 -7760 10580
rect -8230 10514 -8206 10566
rect -8154 10514 -7760 10566
rect -8230 10500 -7760 10514
rect -8810 10200 -8670 10204
rect -8806 10188 -8674 10200
rect -7780 9760 -7640 9920
rect -2992 9258 -2808 9286
rect -2992 9142 -2958 9258
rect -2842 9142 -2808 9258
rect -8630 9106 -8550 9120
rect -2992 9114 -2808 9142
rect -8630 9054 -8616 9106
rect -8564 9054 -8550 9106
rect -8630 9040 -8550 9054
rect -8850 8816 -8770 8820
rect -8850 8810 -8836 8816
rect -13422 8764 -8836 8810
rect -8784 8764 -8770 8816
rect -10600 8760 -10540 8764
rect -8850 8760 -8770 8764
rect -7950 8816 -7870 8820
rect -7950 8764 -7936 8816
rect -7884 8764 -7870 8816
rect -7950 8760 -7870 8764
rect -8700 8200 -4700 8400
rect -10090 7856 -9100 7860
rect -10090 7804 -10076 7856
rect -10024 7804 -9100 7856
rect -10090 7800 -9100 7804
rect -9200 5800 -9100 7800
rect -8710 6076 -8590 6100
rect -8710 6024 -8676 6076
rect -8624 6024 -8590 6076
rect -8710 6000 -8590 6024
rect -13300 5700 -9100 5800
rect -13300 5020 -13200 5700
rect -9200 -100 -9100 5700
rect -4900 4000 -4700 8200
rect -4900 3800 -700 4000
rect 4648 338 5052 366
rect 4648 222 4664 338
rect 5036 222 5052 338
rect 4648 194 5052 222
rect -13300 -200 -9100 -100
rect -13300 -900 -13200 -200
rect -9200 -3200 -9100 -200
rect 6060 -1220 6880 -1160
rect -1566 -2400 -1434 -2388
rect -1570 -2422 -1430 -2400
rect -1570 -2538 -1558 -2422
rect -1442 -2538 -1430 -2422
rect -1570 -2560 -1430 -2538
rect -1566 -2572 -1434 -2560
rect -1770 -2942 -1650 -2940
rect -1770 -2994 -1736 -2942
rect -1684 -2994 -1650 -2942
rect -1770 -3006 -1650 -2994
rect -1770 -3058 -1736 -3006
rect -1684 -3058 -1650 -3006
rect -1770 -3060 -1650 -3058
rect 6060 -3540 6140 -1220
rect 9608 -2842 9932 -2834
rect 9608 -2847 9648 -2842
rect 9892 -2847 9932 -2842
rect 9608 -2953 9645 -2847
rect 9895 -2953 9932 -2847
rect 9608 -2958 9648 -2953
rect 9892 -2958 9932 -2953
rect 8110 -2984 8210 -2960
rect 9608 -2966 9932 -2958
rect 33488 -2842 33812 -2834
rect 33488 -2847 33528 -2842
rect 33772 -2847 33812 -2842
rect 33488 -2953 33525 -2847
rect 33775 -2953 33812 -2847
rect 33488 -2958 33528 -2953
rect 33772 -2958 33812 -2953
rect 33488 -2966 33812 -2958
rect 61788 -2842 62112 -2834
rect 61788 -2847 61828 -2842
rect 62072 -2847 62112 -2842
rect 61788 -2953 61825 -2847
rect 62075 -2953 62112 -2847
rect 61788 -2958 61828 -2953
rect 62072 -2958 62112 -2953
rect 61788 -2966 62112 -2958
rect 8110 -3036 8134 -2984
rect 8186 -3036 8210 -2984
rect 8110 -3060 8210 -3036
rect -14180 -3580 -13640 -3540
rect -14180 -3760 -14118 -3580
rect -13682 -3760 -13640 -3580
rect 6050 -3542 6150 -3540
rect 6050 -3594 6074 -3542
rect 6126 -3594 6150 -3542
rect 6050 -3606 6150 -3594
rect 6050 -3658 6074 -3606
rect 6126 -3658 6150 -3606
rect 6050 -3660 6150 -3658
rect 6600 -3542 7600 -3500
rect 6600 -3594 6654 -3542
rect 6706 -3594 7600 -3542
rect 6600 -3606 7600 -3594
rect 6600 -3658 6654 -3606
rect 6706 -3658 7600 -3606
rect 6060 -3700 6140 -3660
rect 6600 -3700 7600 -3658
rect -14180 -3800 -13640 -3760
rect -11660 -3832 7040 -3800
rect -11660 -3884 6954 -3832
rect 7006 -3884 7040 -3832
rect -11660 -3936 -11476 -3884
rect -11424 -3896 7040 -3884
rect -11424 -3936 6954 -3896
rect -11660 -3948 6954 -3936
rect 7006 -3948 7040 -3896
rect -11660 -4000 7040 -3948
rect 6800 -4500 7040 -4000
rect 6800 -4700 7800 -4500
rect -14200 -9222 -13640 -9020
rect -14200 -9978 -14086 -9222
rect -13714 -9978 -13640 -9222
rect -14200 -10160 -13640 -9978
rect 9590 -10242 9910 -10240
rect 9590 -10358 9628 -10242
rect 9872 -10358 9910 -10242
rect 9590 -10360 9910 -10358
rect 35690 -10242 36006 -10240
rect 35690 -10358 35726 -10242
rect 35970 -10358 36006 -10242
rect 35690 -10360 36006 -10358
rect 61790 -10242 62110 -10240
rect 61790 -10358 61828 -10242
rect 62072 -10358 62110 -10242
rect 61790 -10360 62110 -10358
<< via1 >>
rect -10876 11217 -10824 11230
rect -10876 11183 -10867 11217
rect -10867 11183 -10833 11217
rect -10833 11183 -10824 11217
rect -10876 11178 -10824 11183
rect -10876 11145 -10824 11166
rect -10876 11114 -10867 11145
rect -10867 11114 -10833 11145
rect -10833 11114 -10824 11145
rect 1224 11124 1276 11176
rect -10876 11073 -10824 11102
rect -10876 11050 -10867 11073
rect -10867 11050 -10833 11073
rect -10833 11050 -10824 11073
rect -7736 11054 -7684 11106
rect -10876 11001 -10824 11038
rect -10876 10986 -10867 11001
rect -10867 10986 -10833 11001
rect -10833 10986 -10824 11001
rect -10876 10967 -10867 10974
rect -10867 10967 -10833 10974
rect -10833 10967 -10824 10974
rect -10876 10929 -10824 10967
rect -10876 10922 -10867 10929
rect -10867 10922 -10833 10929
rect -10833 10922 -10824 10929
rect -10876 10895 -10867 10910
rect -10867 10895 -10833 10910
rect -10833 10895 -10824 10910
rect -10876 10858 -10824 10895
rect -10876 10823 -10867 10846
rect -10867 10823 -10833 10846
rect -10833 10823 -10824 10846
rect -10876 10794 -10824 10823
rect -10876 10751 -10867 10782
rect -10867 10751 -10833 10782
rect -10833 10751 -10824 10782
rect -10876 10730 -10824 10751
rect -10876 10713 -10824 10718
rect -10876 10679 -10867 10713
rect -10867 10679 -10833 10713
rect -10833 10679 -10824 10713
rect -10876 10666 -10824 10679
rect -10876 10641 -10824 10654
rect -10876 10607 -10867 10641
rect -10867 10607 -10833 10641
rect -10833 10607 -10824 10641
rect -10876 10602 -10824 10607
rect -10876 10569 -10824 10590
rect -10876 10538 -10867 10569
rect -10867 10538 -10833 10569
rect -10833 10538 -10824 10569
rect -10876 10497 -10824 10526
rect -10876 10474 -10867 10497
rect -10867 10474 -10833 10497
rect -10833 10474 -10824 10497
rect -10876 10425 -10824 10462
rect -10876 10410 -10867 10425
rect -10867 10410 -10833 10425
rect -10833 10410 -10824 10425
rect -10876 10391 -10867 10398
rect -10867 10391 -10833 10398
rect -10833 10391 -10824 10398
rect -10876 10353 -10824 10391
rect -10876 10346 -10867 10353
rect -10867 10346 -10833 10353
rect -10833 10346 -10824 10353
rect -10876 10319 -10867 10334
rect -10867 10319 -10833 10334
rect -10833 10319 -10824 10334
rect -10876 10282 -10824 10319
rect -10876 10247 -10867 10270
rect -10867 10247 -10833 10270
rect -10833 10247 -10824 10270
rect -10876 10218 -10824 10247
rect -10876 10175 -10867 10206
rect -10867 10175 -10833 10206
rect -10833 10175 -10824 10206
rect -10876 10154 -10824 10175
rect -10876 10137 -10824 10142
rect -10876 10103 -10867 10137
rect -10867 10103 -10833 10137
rect -10833 10103 -10824 10137
rect -10876 10090 -10824 10103
rect -8798 10551 -8682 10576
rect -8798 10229 -8793 10551
rect -8793 10229 -8687 10551
rect -8687 10229 -8682 10551
rect -8798 10204 -8682 10229
rect -8206 10514 -8154 10566
rect -2958 9253 -2842 9258
rect -2958 9147 -2953 9253
rect -2953 9147 -2847 9253
rect -2847 9147 -2842 9253
rect -2958 9142 -2842 9147
rect -8616 9054 -8564 9106
rect -8836 8764 -8784 8816
rect -7936 8764 -7884 8816
rect -10076 7804 -10024 7856
rect -8676 6024 -8624 6076
rect 4664 333 5036 338
rect 4664 227 4689 333
rect 4689 227 5011 333
rect 5011 227 5036 333
rect 4664 222 5036 227
rect -1558 -2427 -1442 -2422
rect -1558 -2533 -1553 -2427
rect -1553 -2533 -1447 -2427
rect -1447 -2533 -1442 -2427
rect -1558 -2538 -1442 -2533
rect -1736 -2994 -1684 -2942
rect -1736 -3058 -1684 -3006
rect 9648 -2847 9892 -2842
rect 9648 -2953 9892 -2847
rect 9648 -2958 9892 -2953
rect 33528 -2847 33772 -2842
rect 33528 -2953 33772 -2847
rect 33528 -2958 33772 -2953
rect 61828 -2847 62072 -2842
rect 61828 -2953 62072 -2847
rect 61828 -2958 62072 -2953
rect 8134 -3036 8186 -2984
rect -14118 -3760 -13682 -3580
rect 6074 -3594 6126 -3542
rect 6074 -3658 6126 -3606
rect 6654 -3594 6706 -3542
rect 6654 -3658 6706 -3606
rect 6954 -3884 7006 -3832
rect -11476 -3936 -11424 -3884
rect 6954 -3948 7006 -3896
rect -14086 -9978 -13714 -9222
rect 9628 -10358 9872 -10242
rect 35726 -10358 35970 -10242
rect 61828 -10358 62072 -10242
<< metal2 >>
rect -10900 11248 -10800 11270
rect -10900 11192 -10878 11248
rect -10822 11246 -10800 11248
rect -10822 11192 -10642 11246
rect -10900 11178 -10876 11192
rect -10824 11186 -10642 11192
rect -10824 11178 -10800 11186
rect -10900 11168 -10800 11178
rect -10900 11112 -10878 11168
rect -10822 11112 -10800 11168
rect -7900 11140 -7700 12500
rect 1160 11176 1380 11220
rect -10900 11102 -10800 11112
rect -10900 11088 -10876 11102
rect -10824 11088 -10800 11102
rect -10900 11032 -10878 11088
rect -10822 11032 -10800 11088
rect -10900 11008 -10876 11032
rect -10824 11008 -10800 11032
rect -8940 11106 -7680 11140
rect -8940 11054 -7736 11106
rect -7684 11054 -7680 11106
rect -8940 11020 -7680 11054
rect 1160 11124 1224 11176
rect 1276 11124 1380 11176
rect -10900 10952 -10878 11008
rect -10822 10952 -10800 11008
rect -10900 10928 -10876 10952
rect -10824 10928 -10800 10952
rect -10900 10872 -10878 10928
rect -10822 10886 -10800 10928
rect -10822 10872 -10648 10886
rect -10900 10858 -10876 10872
rect -10824 10858 -10648 10872
rect -10900 10848 -10648 10858
rect -10900 10792 -10878 10848
rect -10822 10826 -10648 10848
rect -8480 10848 -8400 10870
rect -10822 10792 -10800 10826
rect -10900 10782 -10800 10792
rect -10900 10768 -10876 10782
rect -10824 10768 -10800 10782
rect -10900 10712 -10878 10768
rect -10822 10712 -10800 10768
rect -10900 10688 -10876 10712
rect -10824 10688 -10800 10712
rect -10900 10632 -10878 10688
rect -10822 10632 -10800 10688
rect -10900 10608 -10876 10632
rect -10824 10608 -10800 10632
rect -10900 10552 -10878 10608
rect -10822 10552 -10800 10608
rect -8480 10792 -8468 10848
rect -8412 10792 -8400 10848
rect -10900 10538 -10876 10552
rect -10824 10538 -10800 10552
rect -10900 10528 -10800 10538
rect -10900 10472 -10878 10528
rect -10822 10506 -10800 10528
rect -8800 10578 -8680 10590
rect -8800 10576 -8768 10578
rect -8712 10576 -8680 10578
rect -10822 10472 -10656 10506
rect -10900 10462 -10656 10472
rect -10900 10448 -10876 10462
rect -10824 10448 -10656 10462
rect -10900 10392 -10878 10448
rect -10822 10446 -10656 10448
rect -10822 10392 -10800 10446
rect -10900 10368 -10876 10392
rect -10824 10368 -10800 10392
rect -10900 10312 -10878 10368
rect -10822 10312 -10800 10368
rect -10900 10288 -10876 10312
rect -10824 10288 -10800 10312
rect -10900 10232 -10878 10288
rect -10822 10232 -10800 10288
rect -10900 10218 -10876 10232
rect -10824 10218 -10800 10232
rect -10900 10208 -10800 10218
rect -10900 10152 -10878 10208
rect -10822 10152 -10800 10208
rect -8800 10204 -8798 10576
rect -8682 10204 -8680 10576
rect -8800 10202 -8768 10204
rect -8712 10202 -8680 10204
rect -8800 10190 -8680 10202
rect -10900 10146 -10800 10152
rect -10900 10142 -10650 10146
rect -10900 10128 -10876 10142
rect -10824 10128 -10650 10142
rect -10900 10072 -10878 10128
rect -10822 10086 -10650 10128
rect -10822 10072 -10800 10086
rect -10900 9680 -10800 10072
rect -9100 9778 -9000 10000
rect -9100 9722 -9078 9778
rect -9022 9722 -9000 9778
rect -9100 9700 -9000 9722
rect -10900 9620 -10620 9680
rect -10900 9320 -10800 9620
rect -8660 9520 -8600 9530
rect -9440 9518 -8600 9520
rect -9440 9462 -8658 9518
rect -8602 9462 -8600 9518
rect -9440 9460 -8600 9462
rect -8660 9450 -8600 9460
rect -10900 9260 -10620 9320
rect -10900 9240 -10800 9260
rect -14160 8460 -13540 8520
rect -14160 5760 -14100 8460
rect -11260 7680 -11180 8700
rect -10080 7856 -10020 9160
rect -8620 9120 -8560 9130
rect -8480 9120 -8400 10792
rect -8220 10568 -8140 10590
rect -8220 10512 -8208 10568
rect -8152 10512 -8140 10568
rect -8220 10490 -8140 10512
rect -8620 9106 -8400 9120
rect -2980 9268 -2820 9290
rect -2980 9132 -2968 9268
rect -2832 9132 -2820 9268
rect -2980 9110 -2820 9132
rect -8620 9054 -8616 9106
rect -8564 9054 -8400 9106
rect -8620 9040 -8400 9054
rect -8620 9030 -8560 9040
rect -8860 8818 -8760 8850
rect -8860 8762 -8838 8818
rect -8782 8762 -8760 8818
rect -8860 8730 -8760 8762
rect -8216 8840 -8114 8940
rect -8216 8818 -7880 8840
rect -8216 8762 -8198 8818
rect -8142 8816 -7880 8818
rect -8142 8764 -7936 8816
rect -7884 8764 -7880 8816
rect 1160 8800 1380 11124
rect -8142 8762 -7880 8764
rect -8216 8740 -7880 8762
rect -10080 7804 -10076 7856
rect -10024 7804 -10020 7856
rect -10080 7790 -10020 7804
rect -11260 7620 -9480 7680
rect -9540 6100 -9480 7620
rect -8216 6980 -8114 8740
rect 1200 8700 1300 8800
rect -8700 6100 -8600 6110
rect -9540 6076 -8600 6100
rect -9540 6024 -8676 6076
rect -8624 6024 -8600 6076
rect -9540 6000 -8600 6024
rect -11600 5760 -11540 5770
rect -14160 5758 -11540 5760
rect -14160 5702 -11598 5758
rect -11542 5702 -11540 5758
rect -14160 5700 -11540 5702
rect -11600 5690 -11540 5700
rect -11460 5760 -11400 5770
rect -9540 5760 -9480 6000
rect -8700 5990 -8600 6000
rect -11460 5758 -9480 5760
rect -11460 5702 -11458 5758
rect -11402 5702 -9480 5758
rect -11460 5700 -9480 5702
rect -11460 5690 -11400 5700
rect -11460 5118 -11400 5130
rect -11460 5062 -11458 5118
rect -11402 5062 -11400 5118
rect -11460 4280 -11400 5062
rect 6400 4400 28300 4600
rect -11520 4240 -11400 4280
rect -11620 4098 -11500 4126
rect -11620 4042 -11598 4098
rect -11542 4042 -11500 4098
rect -11620 4000 -11500 4042
rect -11280 3178 -11220 3190
rect -11280 3122 -11278 3178
rect -11222 3122 -11220 3178
rect -11280 2500 -11220 3122
rect -11280 2300 1300 2500
rect 1060 1820 1300 2300
rect 4660 348 5040 370
rect 4660 212 4662 348
rect 5038 212 5040 348
rect 6420 308 6600 4400
rect 28000 4300 28300 4400
rect 27200 4100 29100 4300
rect 29400 4228 31300 4300
rect 29400 4172 30242 4228
rect 30298 4172 30322 4228
rect 30378 4172 30402 4228
rect 30458 4172 31300 4228
rect 29400 4100 31300 4172
rect 31600 4228 33500 4300
rect 31600 4172 32442 4228
rect 32498 4172 32522 4228
rect 32578 4172 32602 4228
rect 32658 4172 33500 4228
rect 31600 4100 33500 4172
rect 33800 4228 35700 4300
rect 33800 4172 34642 4228
rect 34698 4172 34722 4228
rect 34778 4172 34802 4228
rect 34858 4172 35700 4228
rect 33800 4100 35700 4172
rect 36000 4228 37900 4300
rect 36000 4172 36842 4228
rect 36898 4172 36922 4228
rect 36978 4172 37002 4228
rect 37058 4172 37900 4228
rect 36000 4100 37900 4172
rect 38200 4228 40100 4300
rect 38200 4172 39042 4228
rect 39098 4172 39122 4228
rect 39178 4172 39202 4228
rect 39258 4172 40100 4228
rect 38200 4100 40100 4172
rect 40400 4228 42300 4300
rect 40400 4172 41242 4228
rect 41298 4172 41322 4228
rect 41378 4172 41402 4228
rect 41458 4172 42300 4228
rect 40400 4100 42300 4172
rect 42600 4228 44500 4300
rect 42600 4172 43442 4228
rect 43498 4172 43522 4228
rect 43578 4172 43602 4228
rect 43658 4172 44500 4228
rect 42600 4100 44500 4172
rect 6420 252 6482 308
rect 6538 252 6600 308
rect 6420 240 6600 252
rect 6480 230 6540 240
rect 4660 190 5040 212
rect 6460 -840 6540 -830
rect 6460 -862 6560 -840
rect 6460 -918 6472 -862
rect 6528 -918 6560 -862
rect 6460 -960 6560 -918
rect 6900 -1472 7060 -1440
rect 6900 -1528 6952 -1472
rect 7008 -1528 7060 -1472
rect 6900 -1540 7060 -1528
rect 6920 -1550 7040 -1540
rect -11540 -1622 -11420 -1600
rect -11540 -1678 -11508 -1622
rect -11452 -1678 -11420 -1622
rect -11540 -1700 -11420 -1678
rect -11880 -1812 -11780 -1790
rect -11880 -1868 -11858 -1812
rect -11802 -1868 -11780 -1812
rect -11880 -1890 -11780 -1868
rect -1560 -2412 -1440 -2390
rect -1560 -2422 -1528 -2412
rect -1472 -2422 -1440 -2412
rect -1560 -2538 -1558 -2422
rect -1442 -2538 -1440 -2422
rect -1560 -2548 -1528 -2538
rect -1472 -2548 -1440 -2538
rect -1560 -2570 -1440 -2548
rect 28000 -2812 28300 -2600
rect 9620 -2842 9920 -2830
rect 9620 -2872 9648 -2842
rect 9892 -2872 9920 -2842
rect -1800 -2942 6720 -2900
rect 9620 -2928 9622 -2872
rect 9918 -2928 9920 -2872
rect 28000 -2868 28042 -2812
rect 28098 -2868 28122 -2812
rect 28178 -2868 28202 -2812
rect 28258 -2868 28300 -2812
rect 28000 -2900 28300 -2868
rect 30200 -2812 30500 -2600
rect 30200 -2868 30242 -2812
rect 30298 -2868 30322 -2812
rect 30378 -2868 30402 -2812
rect 30458 -2868 30500 -2812
rect 30200 -2900 30500 -2868
rect 32400 -2812 32700 -2600
rect 32400 -2868 32442 -2812
rect 32498 -2868 32522 -2812
rect 32578 -2868 32602 -2812
rect 32658 -2868 32700 -2812
rect 34600 -2812 34900 -2600
rect 32400 -2900 32700 -2868
rect 33500 -2842 33800 -2830
rect 33500 -2872 33528 -2842
rect 33772 -2872 33800 -2842
rect -1800 -2994 -1736 -2942
rect -1684 -2994 6720 -2942
rect -5600 -3500 -5400 -3000
rect -1800 -3006 6720 -2994
rect -1800 -3058 -1736 -3006
rect -1684 -3058 6720 -3006
rect -1800 -3100 6720 -3058
rect 6920 -2982 8240 -2940
rect 9620 -2958 9648 -2928
rect 9892 -2958 9920 -2928
rect 9620 -2970 9920 -2958
rect 33500 -2928 33502 -2872
rect 33798 -2928 33800 -2872
rect 34600 -2868 34642 -2812
rect 34698 -2868 34722 -2812
rect 34778 -2868 34802 -2812
rect 34858 -2868 34900 -2812
rect 34600 -2900 34900 -2868
rect 36800 -2812 37100 -2600
rect 36800 -2868 36842 -2812
rect 36898 -2868 36922 -2812
rect 36978 -2868 37002 -2812
rect 37058 -2868 37100 -2812
rect 36800 -2900 37100 -2868
rect 39000 -2812 39300 -2600
rect 39000 -2868 39042 -2812
rect 39098 -2868 39122 -2812
rect 39178 -2868 39202 -2812
rect 39258 -2868 39300 -2812
rect 39000 -2900 39300 -2868
rect 41200 -2812 41500 -2600
rect 41200 -2868 41242 -2812
rect 41298 -2868 41322 -2812
rect 41378 -2868 41402 -2812
rect 41458 -2868 41500 -2812
rect 41200 -2900 41500 -2868
rect 43400 -2812 43700 -2600
rect 43400 -2868 43442 -2812
rect 43498 -2868 43522 -2812
rect 43578 -2868 43602 -2812
rect 43658 -2868 43700 -2812
rect 43400 -2900 43700 -2868
rect 61800 -2842 62100 -2830
rect 61800 -2872 61828 -2842
rect 62072 -2872 62100 -2842
rect 33500 -2958 33528 -2928
rect 33772 -2958 33800 -2928
rect 33500 -2970 33800 -2958
rect 61800 -2928 61802 -2872
rect 62098 -2928 62100 -2872
rect 61800 -2958 61828 -2928
rect 62072 -2958 62100 -2928
rect 61800 -2970 62100 -2958
rect 6920 -3038 6952 -2982
rect 7008 -2984 8240 -2982
rect 7008 -3036 8134 -2984
rect 8186 -3036 8240 -2984
rect 7008 -3038 8240 -3036
rect 6920 -3080 8240 -3038
rect -5600 -3542 6200 -3500
rect -14140 -3562 -13660 -3550
rect -14140 -3778 -14128 -3562
rect -13672 -3778 -13660 -3562
rect -5600 -3594 6074 -3542
rect 6126 -3594 6200 -3542
rect -5600 -3606 6200 -3594
rect -5600 -3658 6074 -3606
rect 6126 -3658 6200 -3606
rect -5600 -3700 6200 -3658
rect 6600 -3542 6720 -3100
rect 6600 -3594 6654 -3542
rect 6706 -3594 6720 -3542
rect 6600 -3606 6720 -3594
rect 6600 -3658 6654 -3606
rect 6706 -3658 6720 -3606
rect 6600 -3680 6720 -3658
rect -14140 -3790 -13660 -3778
rect 6940 -3822 7020 -3790
rect -11500 -3882 -11400 -3850
rect -11500 -3938 -11478 -3882
rect -11422 -3938 -11400 -3882
rect -11500 -3970 -11400 -3938
rect 6940 -3878 6952 -3822
rect 7008 -3878 7020 -3822
rect 6940 -3884 6954 -3878
rect 7006 -3884 7020 -3878
rect 6940 -3896 7020 -3884
rect 6940 -3902 6954 -3896
rect 7006 -3902 7020 -3896
rect 6940 -3958 6952 -3902
rect 7008 -3958 7020 -3902
rect 6940 -3990 7020 -3958
rect -14100 -9212 -13700 -9190
rect -14100 -9988 -14088 -9212
rect -13712 -9988 -13700 -9212
rect -14100 -10010 -13700 -9988
rect 9600 -10242 9900 -10230
rect 9600 -10272 9628 -10242
rect 9872 -10272 9900 -10242
rect 9600 -10328 9602 -10272
rect 9898 -10328 9900 -10272
rect 9600 -10358 9628 -10328
rect 9872 -10358 9900 -10328
rect 9600 -10370 9900 -10358
rect 35700 -10242 35996 -10230
rect 35700 -10272 35726 -10242
rect 35970 -10272 35996 -10242
rect 35700 -10358 35726 -10328
rect 35970 -10358 35996 -10328
rect 35700 -10370 35996 -10358
rect 61800 -10242 62100 -10230
rect 61800 -10272 61828 -10242
rect 62072 -10272 62100 -10242
rect 61800 -10328 61802 -10272
rect 62098 -10328 62100 -10272
rect 61800 -10358 61828 -10328
rect 62072 -10358 62100 -10328
rect 61800 -10370 62100 -10358
<< via2 >>
rect -10878 11230 -10822 11248
rect -10878 11192 -10876 11230
rect -10876 11192 -10824 11230
rect -10824 11192 -10822 11230
rect -10878 11166 -10822 11168
rect -10878 11114 -10876 11166
rect -10876 11114 -10824 11166
rect -10824 11114 -10822 11166
rect -10878 11112 -10822 11114
rect -10878 11050 -10876 11088
rect -10876 11050 -10824 11088
rect -10824 11050 -10822 11088
rect -10878 11038 -10822 11050
rect -10878 11032 -10876 11038
rect -10876 11032 -10824 11038
rect -10824 11032 -10822 11038
rect -10878 10986 -10876 11008
rect -10876 10986 -10824 11008
rect -10824 10986 -10822 11008
rect -10878 10974 -10822 10986
rect -10878 10952 -10876 10974
rect -10876 10952 -10824 10974
rect -10824 10952 -10822 10974
rect -10878 10922 -10876 10928
rect -10876 10922 -10824 10928
rect -10824 10922 -10822 10928
rect -10878 10910 -10822 10922
rect -10878 10872 -10876 10910
rect -10876 10872 -10824 10910
rect -10824 10872 -10822 10910
rect -10878 10846 -10822 10848
rect -10878 10794 -10876 10846
rect -10876 10794 -10824 10846
rect -10824 10794 -10822 10846
rect -10878 10792 -10822 10794
rect -10878 10730 -10876 10768
rect -10876 10730 -10824 10768
rect -10824 10730 -10822 10768
rect -10878 10718 -10822 10730
rect -10878 10712 -10876 10718
rect -10876 10712 -10824 10718
rect -10824 10712 -10822 10718
rect -10878 10666 -10876 10688
rect -10876 10666 -10824 10688
rect -10824 10666 -10822 10688
rect -10878 10654 -10822 10666
rect -10878 10632 -10876 10654
rect -10876 10632 -10824 10654
rect -10824 10632 -10822 10654
rect -10878 10602 -10876 10608
rect -10876 10602 -10824 10608
rect -10824 10602 -10822 10608
rect -10878 10590 -10822 10602
rect -10878 10552 -10876 10590
rect -10876 10552 -10824 10590
rect -10824 10552 -10822 10590
rect -8468 10792 -8412 10848
rect -10878 10526 -10822 10528
rect -10878 10474 -10876 10526
rect -10876 10474 -10824 10526
rect -10824 10474 -10822 10526
rect -8768 10576 -8712 10578
rect -10878 10472 -10822 10474
rect -10878 10410 -10876 10448
rect -10876 10410 -10824 10448
rect -10824 10410 -10822 10448
rect -10878 10398 -10822 10410
rect -10878 10392 -10876 10398
rect -10876 10392 -10824 10398
rect -10824 10392 -10822 10398
rect -10878 10346 -10876 10368
rect -10876 10346 -10824 10368
rect -10824 10346 -10822 10368
rect -10878 10334 -10822 10346
rect -10878 10312 -10876 10334
rect -10876 10312 -10824 10334
rect -10824 10312 -10822 10334
rect -10878 10282 -10876 10288
rect -10876 10282 -10824 10288
rect -10824 10282 -10822 10288
rect -10878 10270 -10822 10282
rect -10878 10232 -10876 10270
rect -10876 10232 -10824 10270
rect -10824 10232 -10822 10270
rect -10878 10206 -10822 10208
rect -10878 10154 -10876 10206
rect -10876 10154 -10824 10206
rect -10824 10154 -10822 10206
rect -10878 10152 -10822 10154
rect -8768 10522 -8712 10576
rect -8768 10442 -8712 10498
rect -8768 10362 -8712 10418
rect -8768 10282 -8712 10338
rect -8768 10204 -8712 10258
rect -8768 10202 -8712 10204
rect -10878 10090 -10876 10128
rect -10876 10090 -10824 10128
rect -10824 10090 -10822 10128
rect -10878 10072 -10822 10090
rect -9078 9722 -9022 9778
rect -8658 9462 -8602 9518
rect -8208 10566 -8152 10568
rect -8208 10514 -8206 10566
rect -8206 10514 -8154 10566
rect -8154 10514 -8152 10566
rect -8208 10512 -8152 10514
rect -2968 9258 -2832 9268
rect -2968 9142 -2958 9258
rect -2958 9142 -2842 9258
rect -2842 9142 -2832 9258
rect -2968 9132 -2832 9142
rect -8838 8816 -8782 8818
rect -8838 8764 -8836 8816
rect -8836 8764 -8784 8816
rect -8784 8764 -8782 8816
rect -8838 8762 -8782 8764
rect -8198 8762 -8142 8818
rect -11598 5702 -11542 5758
rect -11458 5702 -11402 5758
rect -11458 5062 -11402 5118
rect -11598 4042 -11542 4098
rect -11278 3122 -11222 3178
rect 4662 338 5038 348
rect 4662 222 4664 338
rect 4664 222 5036 338
rect 5036 222 5038 338
rect 4662 212 5038 222
rect 30242 4172 30298 4228
rect 30322 4172 30378 4228
rect 30402 4172 30458 4228
rect 32442 4172 32498 4228
rect 32522 4172 32578 4228
rect 32602 4172 32658 4228
rect 34642 4172 34698 4228
rect 34722 4172 34778 4228
rect 34802 4172 34858 4228
rect 36842 4172 36898 4228
rect 36922 4172 36978 4228
rect 37002 4172 37058 4228
rect 39042 4172 39098 4228
rect 39122 4172 39178 4228
rect 39202 4172 39258 4228
rect 41242 4172 41298 4228
rect 41322 4172 41378 4228
rect 41402 4172 41458 4228
rect 43442 4172 43498 4228
rect 43522 4172 43578 4228
rect 43602 4172 43658 4228
rect 6482 252 6538 308
rect 6472 -918 6528 -862
rect 6952 -1528 7008 -1472
rect -11508 -1678 -11452 -1622
rect -11858 -1868 -11802 -1812
rect -1528 -2422 -1472 -2412
rect -1528 -2468 -1472 -2422
rect -1528 -2538 -1472 -2492
rect -1528 -2548 -1472 -2538
rect 9622 -2928 9648 -2872
rect 9648 -2928 9678 -2872
rect 9702 -2928 9758 -2872
rect 9782 -2928 9838 -2872
rect 9862 -2928 9892 -2872
rect 9892 -2928 9918 -2872
rect 28042 -2868 28098 -2812
rect 28122 -2868 28178 -2812
rect 28202 -2868 28258 -2812
rect 30242 -2868 30298 -2812
rect 30322 -2868 30378 -2812
rect 30402 -2868 30458 -2812
rect 32442 -2868 32498 -2812
rect 32522 -2868 32578 -2812
rect 32602 -2868 32658 -2812
rect 33502 -2928 33528 -2872
rect 33528 -2928 33558 -2872
rect 33582 -2928 33638 -2872
rect 33662 -2928 33718 -2872
rect 33742 -2928 33772 -2872
rect 33772 -2928 33798 -2872
rect 34642 -2868 34698 -2812
rect 34722 -2868 34778 -2812
rect 34802 -2868 34858 -2812
rect 36842 -2868 36898 -2812
rect 36922 -2868 36978 -2812
rect 37002 -2868 37058 -2812
rect 39042 -2868 39098 -2812
rect 39122 -2868 39178 -2812
rect 39202 -2868 39258 -2812
rect 41242 -2868 41298 -2812
rect 41322 -2868 41378 -2812
rect 41402 -2868 41458 -2812
rect 43442 -2868 43498 -2812
rect 43522 -2868 43578 -2812
rect 43602 -2868 43658 -2812
rect 61802 -2928 61828 -2872
rect 61828 -2928 61858 -2872
rect 61882 -2928 61938 -2872
rect 61962 -2928 62018 -2872
rect 62042 -2928 62072 -2872
rect 62072 -2928 62098 -2872
rect 6952 -3038 7008 -2982
rect -14128 -3580 -13672 -3562
rect -14128 -3760 -14118 -3580
rect -14118 -3760 -13682 -3580
rect -13682 -3760 -13672 -3580
rect -14128 -3778 -13672 -3760
rect -11478 -3884 -11422 -3882
rect -11478 -3936 -11476 -3884
rect -11476 -3936 -11424 -3884
rect -11424 -3936 -11422 -3884
rect -11478 -3938 -11422 -3936
rect 6952 -3832 7008 -3822
rect 6952 -3878 6954 -3832
rect 6954 -3878 7006 -3832
rect 7006 -3878 7008 -3832
rect 6952 -3948 6954 -3902
rect 6954 -3948 7006 -3902
rect 7006 -3948 7008 -3902
rect 6952 -3958 7008 -3948
rect -14088 -9222 -13712 -9212
rect -14088 -9978 -14086 -9222
rect -14086 -9978 -13714 -9222
rect -13714 -9978 -13712 -9222
rect -14088 -9988 -13712 -9978
rect 9602 -10328 9628 -10272
rect 9628 -10328 9658 -10272
rect 9682 -10328 9738 -10272
rect 9762 -10328 9818 -10272
rect 9842 -10328 9872 -10272
rect 9872 -10328 9898 -10272
rect 35700 -10328 35726 -10272
rect 35726 -10328 35756 -10272
rect 35780 -10328 35836 -10272
rect 35860 -10328 35916 -10272
rect 35940 -10328 35970 -10272
rect 35970 -10328 35996 -10272
rect 61802 -10328 61828 -10272
rect 61828 -10328 61858 -10272
rect 61882 -10328 61938 -10272
rect 61962 -10328 62018 -10272
rect 62042 -10328 62072 -10272
rect 62072 -10328 62098 -10272
<< metal3 >>
rect -10910 11252 -10790 11265
rect -10910 11188 -10882 11252
rect -10818 11188 -10790 11252
rect -10910 11172 -10790 11188
rect -10910 11108 -10882 11172
rect -10818 11108 -10790 11172
rect -10910 11092 -10790 11108
rect -10910 11028 -10882 11092
rect -10818 11028 -10790 11092
rect -10910 11012 -10790 11028
rect -10910 10948 -10882 11012
rect -10818 10948 -10790 11012
rect -10910 10932 -10790 10948
rect -10910 10868 -10882 10932
rect -10818 10868 -10790 10932
rect -10910 10852 -10790 10868
rect -10910 10788 -10882 10852
rect -10818 10788 -10790 10852
rect -10910 10772 -10790 10788
rect -10910 10708 -10882 10772
rect -10818 10708 -10790 10772
rect -8500 10848 -8380 12540
rect -8500 10792 -8468 10848
rect -8412 10792 -8380 10848
rect -8500 10760 -8380 10792
rect -10910 10692 -10790 10708
rect -10910 10628 -10882 10692
rect -10818 10628 -10790 10692
rect -10910 10612 -10790 10628
rect -10910 10548 -10882 10612
rect -10818 10548 -10790 10612
rect -10910 10532 -10790 10548
rect -10910 10468 -10882 10532
rect -10818 10468 -10790 10532
rect -10910 10452 -10790 10468
rect -10910 10388 -10882 10452
rect -10818 10388 -10790 10452
rect -10910 10372 -10790 10388
rect -10910 10308 -10882 10372
rect -10818 10308 -10790 10372
rect -10910 10292 -10790 10308
rect -10910 10228 -10882 10292
rect -10818 10228 -10790 10292
rect -10910 10212 -10790 10228
rect -10910 10148 -10882 10212
rect -10818 10148 -10790 10212
rect -8810 10578 -8670 10585
rect -8810 10542 -8768 10578
rect -8712 10542 -8670 10578
rect -8810 10478 -8772 10542
rect -8708 10478 -8670 10542
rect -8230 10568 -8130 10585
rect -8230 10512 -8208 10568
rect -8152 10512 -8130 10568
rect -8230 10495 -8130 10512
rect -8810 10462 -8768 10478
rect -8712 10462 -8670 10478
rect -8810 10398 -8772 10462
rect -8708 10398 -8670 10462
rect -8810 10382 -8768 10398
rect -8712 10382 -8670 10398
rect -8810 10318 -8772 10382
rect -8708 10318 -8670 10382
rect -8810 10302 -8768 10318
rect -8712 10302 -8670 10318
rect -8810 10238 -8772 10302
rect -8708 10238 -8670 10302
rect -8810 10202 -8768 10238
rect -8712 10202 -8670 10238
rect -8810 10195 -8670 10202
rect -10910 10132 -10790 10148
rect -10910 10068 -10882 10132
rect -10818 10068 -10790 10132
rect -10910 10055 -10790 10068
rect -9100 9778 -9000 9800
rect -14190 9726 -14050 9760
rect -10910 9726 -10790 9740
rect -14200 9722 -13460 9726
rect -14200 9666 -14152 9722
rect -14190 9658 -14152 9666
rect -14088 9666 -13460 9722
rect -11340 9722 -10790 9726
rect -11340 9666 -10882 9722
rect -14088 9658 -14050 9666
rect -14190 9620 -14050 9658
rect -10910 9658 -10882 9666
rect -10818 9658 -10790 9722
rect -10910 9640 -10790 9658
rect -9100 9722 -9078 9778
rect -9022 9722 -9000 9778
rect -11610 5758 -11530 5790
rect -11610 5702 -11598 5758
rect -11542 5702 -11530 5758
rect -11610 4098 -11530 5702
rect -11470 5758 -11390 5770
rect -11470 5702 -11458 5758
rect -11402 5702 -11390 5758
rect -11470 5118 -11390 5702
rect -11470 5062 -11458 5118
rect -11402 5062 -11390 5118
rect -11470 5050 -11390 5062
rect -11610 4042 -11598 4098
rect -11542 4042 -11530 4098
rect -11610 3200 -11530 4042
rect -11610 3178 -11200 3200
rect -11610 3122 -11278 3178
rect -11222 3122 -11200 3178
rect -11610 3120 -11200 3122
rect -11290 3115 -11210 3120
rect -9100 2200 -9000 9722
rect -8220 9540 -8140 10495
rect -8680 9518 -8140 9540
rect -8680 9462 -8658 9518
rect -8602 9462 -8140 9518
rect -8680 9440 -8140 9462
rect -2990 9272 -2810 9285
rect -2990 9128 -2972 9272
rect -2828 9128 -2810 9272
rect -2990 9115 -2810 9128
rect -8870 8840 -8750 8845
rect -8870 8818 -8120 8840
rect -8870 8762 -8838 8818
rect -8782 8762 -8198 8818
rect -8142 8762 -8120 8818
rect -8870 8740 -8120 8762
rect -8870 8735 -8750 8740
rect 30200 4228 30500 12600
rect 30200 4172 30242 4228
rect 30298 4172 30322 4228
rect 30378 4172 30402 4228
rect 30458 4172 30500 4228
rect 30200 4100 30500 4172
rect 32400 4228 32700 12600
rect 32400 4172 32442 4228
rect 32498 4172 32522 4228
rect 32578 4172 32602 4228
rect 32658 4172 32700 4228
rect 32400 4100 32700 4172
rect 34600 4228 34900 12600
rect 34600 4172 34642 4228
rect 34698 4172 34722 4228
rect 34778 4172 34802 4228
rect 34858 4172 34900 4228
rect 34600 4100 34900 4172
rect 36800 4228 37100 12600
rect 36800 4172 36842 4228
rect 36898 4172 36922 4228
rect 36978 4172 37002 4228
rect 37058 4172 37100 4228
rect 36800 4100 37100 4172
rect 39000 4228 39300 12600
rect 39000 4172 39042 4228
rect 39098 4172 39122 4228
rect 39178 4172 39202 4228
rect 39258 4172 39300 4228
rect 39000 4100 39300 4172
rect 41200 4228 41500 12600
rect 41200 4172 41242 4228
rect 41298 4172 41322 4228
rect 41378 4172 41402 4228
rect 41458 4172 41500 4228
rect 41200 4100 41500 4172
rect 43400 4228 43700 12600
rect 43400 4172 43442 4228
rect 43498 4172 43522 4228
rect 43578 4172 43602 4228
rect 43658 4172 43700 4228
rect 43400 4100 43700 4172
rect -7040 3212 -6880 4060
rect -7040 3148 -6992 3212
rect -6928 3148 -6880 3212
rect -7040 3132 -6880 3148
rect -7040 3068 -6992 3132
rect -6928 3068 -6880 3132
rect -7040 2200 -6880 3068
rect -11900 2100 -9000 2200
rect -11900 -1795 -11800 2100
rect 4650 352 5050 365
rect 4650 348 4698 352
rect 5002 348 5050 352
rect 4650 212 4662 348
rect 5038 212 5050 348
rect 4650 208 4698 212
rect 5002 208 5050 212
rect 4650 195 5050 208
rect 6460 308 6560 340
rect 6460 252 6482 308
rect 6538 252 6560 308
rect 6460 -835 6560 252
rect 6450 -862 6560 -835
rect 6450 -918 6472 -862
rect 6528 -918 6560 -862
rect 6450 -940 6560 -918
rect 6450 -945 6550 -940
rect 6910 -1472 7050 -1455
rect 6910 -1528 6952 -1472
rect 7008 -1528 7050 -1472
rect 6910 -1545 7050 -1528
rect -11480 -1615 -11420 -1600
rect -11530 -1622 -11420 -1615
rect -11530 -1678 -11508 -1622
rect -11452 -1678 -11420 -1622
rect -11530 -1685 -11420 -1678
rect -11900 -1812 -11770 -1795
rect -11900 -1868 -11858 -1812
rect -11802 -1868 -11770 -1812
rect -11900 -1885 -11770 -1868
rect -11900 -1900 -11800 -1885
rect -14150 -3562 -13650 -3555
rect -14150 -3598 -14128 -3562
rect -13672 -3598 -13650 -3562
rect -14150 -3742 -14132 -3598
rect -13668 -3742 -13650 -3598
rect -14150 -3778 -14128 -3742
rect -13672 -3778 -13650 -3742
rect -14150 -3785 -13650 -3778
rect -11480 -3855 -11420 -1685
rect -1570 -2408 -1430 -2395
rect -1570 -2472 -1532 -2408
rect -1468 -2472 -1430 -2408
rect -1570 -2488 -1430 -2472
rect -1570 -2552 -1532 -2488
rect -1468 -2552 -1430 -2488
rect -1570 -2565 -1430 -2552
rect 6920 -2982 7040 -1545
rect 28030 -2808 28270 -2795
rect 28030 -2812 28078 -2808
rect 28142 -2812 28158 -2808
rect 28222 -2812 28270 -2808
rect 9610 -2868 9930 -2835
rect 9610 -2872 9658 -2868
rect 9722 -2872 9738 -2868
rect 9802 -2872 9818 -2868
rect 9882 -2872 9930 -2868
rect 9610 -2928 9622 -2872
rect 9918 -2928 9930 -2872
rect 28030 -2868 28042 -2812
rect 28258 -2868 28270 -2812
rect 28030 -2872 28078 -2868
rect 28142 -2872 28158 -2868
rect 28222 -2872 28270 -2868
rect 28030 -2885 28270 -2872
rect 30230 -2808 30470 -2795
rect 30230 -2812 30278 -2808
rect 30342 -2812 30358 -2808
rect 30422 -2812 30470 -2808
rect 30230 -2868 30242 -2812
rect 30458 -2868 30470 -2812
rect 30230 -2872 30278 -2868
rect 30342 -2872 30358 -2868
rect 30422 -2872 30470 -2868
rect 30230 -2885 30470 -2872
rect 32430 -2808 32670 -2795
rect 32430 -2812 32478 -2808
rect 32542 -2812 32558 -2808
rect 32622 -2812 32670 -2808
rect 32430 -2868 32442 -2812
rect 32658 -2868 32670 -2812
rect 34630 -2808 34870 -2795
rect 34630 -2812 34678 -2808
rect 34742 -2812 34758 -2808
rect 34822 -2812 34870 -2808
rect 32430 -2872 32478 -2868
rect 32542 -2872 32558 -2868
rect 32622 -2872 32670 -2868
rect 32430 -2885 32670 -2872
rect 33490 -2868 33810 -2835
rect 33490 -2872 33538 -2868
rect 33602 -2872 33618 -2868
rect 33682 -2872 33698 -2868
rect 33762 -2872 33810 -2868
rect 9610 -2932 9658 -2928
rect 9722 -2932 9738 -2928
rect 9802 -2932 9818 -2928
rect 9882 -2932 9930 -2928
rect 9610 -2965 9930 -2932
rect 33490 -2928 33502 -2872
rect 33798 -2928 33810 -2872
rect 34630 -2868 34642 -2812
rect 34858 -2868 34870 -2812
rect 34630 -2872 34678 -2868
rect 34742 -2872 34758 -2868
rect 34822 -2872 34870 -2868
rect 34630 -2885 34870 -2872
rect 36830 -2808 37070 -2795
rect 36830 -2812 36878 -2808
rect 36942 -2812 36958 -2808
rect 37022 -2812 37070 -2808
rect 36830 -2868 36842 -2812
rect 37058 -2868 37070 -2812
rect 36830 -2872 36878 -2868
rect 36942 -2872 36958 -2868
rect 37022 -2872 37070 -2868
rect 36830 -2885 37070 -2872
rect 39030 -2808 39270 -2795
rect 39030 -2812 39078 -2808
rect 39142 -2812 39158 -2808
rect 39222 -2812 39270 -2808
rect 39030 -2868 39042 -2812
rect 39258 -2868 39270 -2812
rect 39030 -2872 39078 -2868
rect 39142 -2872 39158 -2868
rect 39222 -2872 39270 -2868
rect 39030 -2885 39270 -2872
rect 41230 -2808 41470 -2795
rect 41230 -2812 41278 -2808
rect 41342 -2812 41358 -2808
rect 41422 -2812 41470 -2808
rect 41230 -2868 41242 -2812
rect 41458 -2868 41470 -2812
rect 41230 -2872 41278 -2868
rect 41342 -2872 41358 -2868
rect 41422 -2872 41470 -2868
rect 41230 -2885 41470 -2872
rect 43430 -2808 43670 -2795
rect 43430 -2812 43478 -2808
rect 43542 -2812 43558 -2808
rect 43622 -2812 43670 -2808
rect 43430 -2868 43442 -2812
rect 43658 -2868 43670 -2812
rect 43430 -2872 43478 -2868
rect 43542 -2872 43558 -2868
rect 43622 -2872 43670 -2868
rect 43430 -2885 43670 -2872
rect 61790 -2868 62110 -2835
rect 61790 -2872 61838 -2868
rect 61902 -2872 61918 -2868
rect 61982 -2872 61998 -2868
rect 62062 -2872 62110 -2868
rect 33490 -2932 33538 -2928
rect 33602 -2932 33618 -2928
rect 33682 -2932 33698 -2928
rect 33762 -2932 33810 -2928
rect 33490 -2965 33810 -2932
rect 61790 -2928 61802 -2872
rect 62098 -2928 62110 -2872
rect 61790 -2932 61838 -2928
rect 61902 -2932 61918 -2928
rect 61982 -2932 61998 -2928
rect 62062 -2932 62110 -2928
rect 61790 -2965 62110 -2932
rect 6920 -3038 6952 -2982
rect 7008 -3038 7040 -2982
rect 6920 -3822 7040 -3038
rect -11510 -3882 -11390 -3855
rect -11510 -3938 -11478 -3882
rect -11422 -3938 -11390 -3882
rect -11510 -3965 -11390 -3938
rect 6920 -3878 6952 -3822
rect 7008 -3878 7040 -3822
rect 6920 -3902 7040 -3878
rect 6920 -3958 6952 -3902
rect 7008 -3958 7040 -3902
rect 6920 -4000 7040 -3958
rect -14110 -9208 -13690 -9195
rect -14110 -9992 -14092 -9208
rect -13708 -9992 -13690 -9208
rect -14110 -10005 -13690 -9992
rect 9590 -10268 9910 -10235
rect 9590 -10272 9638 -10268
rect 9702 -10272 9718 -10268
rect 9782 -10272 9798 -10268
rect 9862 -10272 9910 -10268
rect 9590 -10328 9602 -10272
rect 9898 -10328 9910 -10272
rect 9590 -10332 9638 -10328
rect 9702 -10332 9718 -10328
rect 9782 -10332 9798 -10328
rect 9862 -10332 9910 -10328
rect 9590 -10365 9910 -10332
rect 35690 -10268 36006 -10235
rect 35690 -10272 35736 -10268
rect 35800 -10272 35816 -10268
rect 35880 -10272 35896 -10268
rect 35960 -10272 36006 -10268
rect 35690 -10328 35700 -10272
rect 35996 -10328 36006 -10272
rect 35690 -10332 35736 -10328
rect 35800 -10332 35816 -10328
rect 35880 -10332 35896 -10328
rect 35960 -10332 36006 -10328
rect 35690 -10365 36006 -10332
rect 61790 -10268 62110 -10235
rect 61790 -10272 61838 -10268
rect 61902 -10272 61918 -10268
rect 61982 -10272 61998 -10268
rect 62062 -10272 62110 -10268
rect 61790 -10328 61802 -10272
rect 62098 -10328 62110 -10272
rect 61790 -10332 61838 -10328
rect 61902 -10332 61918 -10328
rect 61982 -10332 61998 -10328
rect 62062 -10332 62110 -10328
rect 61790 -10365 62110 -10332
<< via3 >>
rect -10882 11248 -10818 11252
rect -10882 11192 -10878 11248
rect -10878 11192 -10822 11248
rect -10822 11192 -10818 11248
rect -10882 11188 -10818 11192
rect -10882 11168 -10818 11172
rect -10882 11112 -10878 11168
rect -10878 11112 -10822 11168
rect -10822 11112 -10818 11168
rect -10882 11108 -10818 11112
rect -10882 11088 -10818 11092
rect -10882 11032 -10878 11088
rect -10878 11032 -10822 11088
rect -10822 11032 -10818 11088
rect -10882 11028 -10818 11032
rect -10882 11008 -10818 11012
rect -10882 10952 -10878 11008
rect -10878 10952 -10822 11008
rect -10822 10952 -10818 11008
rect -10882 10948 -10818 10952
rect -10882 10928 -10818 10932
rect -10882 10872 -10878 10928
rect -10878 10872 -10822 10928
rect -10822 10872 -10818 10928
rect -10882 10868 -10818 10872
rect -10882 10848 -10818 10852
rect -10882 10792 -10878 10848
rect -10878 10792 -10822 10848
rect -10822 10792 -10818 10848
rect -10882 10788 -10818 10792
rect -10882 10768 -10818 10772
rect -10882 10712 -10878 10768
rect -10878 10712 -10822 10768
rect -10822 10712 -10818 10768
rect -10882 10708 -10818 10712
rect -10882 10688 -10818 10692
rect -10882 10632 -10878 10688
rect -10878 10632 -10822 10688
rect -10822 10632 -10818 10688
rect -10882 10628 -10818 10632
rect -10882 10608 -10818 10612
rect -10882 10552 -10878 10608
rect -10878 10552 -10822 10608
rect -10822 10552 -10818 10608
rect -10882 10548 -10818 10552
rect -10882 10528 -10818 10532
rect -10882 10472 -10878 10528
rect -10878 10472 -10822 10528
rect -10822 10472 -10818 10528
rect -10882 10468 -10818 10472
rect -10882 10448 -10818 10452
rect -10882 10392 -10878 10448
rect -10878 10392 -10822 10448
rect -10822 10392 -10818 10448
rect -10882 10388 -10818 10392
rect -10882 10368 -10818 10372
rect -10882 10312 -10878 10368
rect -10878 10312 -10822 10368
rect -10822 10312 -10818 10368
rect -10882 10308 -10818 10312
rect -10882 10288 -10818 10292
rect -10882 10232 -10878 10288
rect -10878 10232 -10822 10288
rect -10822 10232 -10818 10288
rect -10882 10228 -10818 10232
rect -10882 10208 -10818 10212
rect -10882 10152 -10878 10208
rect -10878 10152 -10822 10208
rect -10822 10152 -10818 10208
rect -10882 10148 -10818 10152
rect -8772 10522 -8768 10542
rect -8768 10522 -8712 10542
rect -8712 10522 -8708 10542
rect -8772 10498 -8708 10522
rect -8772 10478 -8768 10498
rect -8768 10478 -8712 10498
rect -8712 10478 -8708 10498
rect -8772 10442 -8768 10462
rect -8768 10442 -8712 10462
rect -8712 10442 -8708 10462
rect -8772 10418 -8708 10442
rect -8772 10398 -8768 10418
rect -8768 10398 -8712 10418
rect -8712 10398 -8708 10418
rect -8772 10362 -8768 10382
rect -8768 10362 -8712 10382
rect -8712 10362 -8708 10382
rect -8772 10338 -8708 10362
rect -8772 10318 -8768 10338
rect -8768 10318 -8712 10338
rect -8712 10318 -8708 10338
rect -8772 10282 -8768 10302
rect -8768 10282 -8712 10302
rect -8712 10282 -8708 10302
rect -8772 10258 -8708 10282
rect -8772 10238 -8768 10258
rect -8768 10238 -8712 10258
rect -8712 10238 -8708 10258
rect -10882 10128 -10818 10132
rect -10882 10072 -10878 10128
rect -10878 10072 -10822 10128
rect -10822 10072 -10818 10128
rect -10882 10068 -10818 10072
rect -14152 9658 -14088 9722
rect -10882 9658 -10818 9722
rect -2972 9268 -2828 9272
rect -2972 9132 -2968 9268
rect -2968 9132 -2832 9268
rect -2832 9132 -2828 9268
rect -2972 9128 -2828 9132
rect -6992 3148 -6928 3212
rect -6992 3068 -6928 3132
rect 4698 348 5002 352
rect 4698 212 5002 348
rect 4698 208 5002 212
rect -14132 -3742 -14128 -3598
rect -14128 -3742 -13672 -3598
rect -13672 -3742 -13668 -3598
rect -1532 -2412 -1468 -2408
rect -1532 -2468 -1528 -2412
rect -1528 -2468 -1472 -2412
rect -1472 -2468 -1468 -2412
rect -1532 -2472 -1468 -2468
rect -1532 -2492 -1468 -2488
rect -1532 -2548 -1528 -2492
rect -1528 -2548 -1472 -2492
rect -1472 -2548 -1468 -2492
rect -1532 -2552 -1468 -2548
rect 28078 -2812 28142 -2808
rect 28158 -2812 28222 -2808
rect 9658 -2872 9722 -2868
rect 9738 -2872 9802 -2868
rect 9818 -2872 9882 -2868
rect 9658 -2928 9678 -2872
rect 9678 -2928 9702 -2872
rect 9702 -2928 9722 -2872
rect 9738 -2928 9758 -2872
rect 9758 -2928 9782 -2872
rect 9782 -2928 9802 -2872
rect 9818 -2928 9838 -2872
rect 9838 -2928 9862 -2872
rect 9862 -2928 9882 -2872
rect 28078 -2868 28098 -2812
rect 28098 -2868 28122 -2812
rect 28122 -2868 28142 -2812
rect 28158 -2868 28178 -2812
rect 28178 -2868 28202 -2812
rect 28202 -2868 28222 -2812
rect 28078 -2872 28142 -2868
rect 28158 -2872 28222 -2868
rect 30278 -2812 30342 -2808
rect 30358 -2812 30422 -2808
rect 30278 -2868 30298 -2812
rect 30298 -2868 30322 -2812
rect 30322 -2868 30342 -2812
rect 30358 -2868 30378 -2812
rect 30378 -2868 30402 -2812
rect 30402 -2868 30422 -2812
rect 30278 -2872 30342 -2868
rect 30358 -2872 30422 -2868
rect 32478 -2812 32542 -2808
rect 32558 -2812 32622 -2808
rect 32478 -2868 32498 -2812
rect 32498 -2868 32522 -2812
rect 32522 -2868 32542 -2812
rect 32558 -2868 32578 -2812
rect 32578 -2868 32602 -2812
rect 32602 -2868 32622 -2812
rect 34678 -2812 34742 -2808
rect 34758 -2812 34822 -2808
rect 32478 -2872 32542 -2868
rect 32558 -2872 32622 -2868
rect 33538 -2872 33602 -2868
rect 33618 -2872 33682 -2868
rect 33698 -2872 33762 -2868
rect 9658 -2932 9722 -2928
rect 9738 -2932 9802 -2928
rect 9818 -2932 9882 -2928
rect 33538 -2928 33558 -2872
rect 33558 -2928 33582 -2872
rect 33582 -2928 33602 -2872
rect 33618 -2928 33638 -2872
rect 33638 -2928 33662 -2872
rect 33662 -2928 33682 -2872
rect 33698 -2928 33718 -2872
rect 33718 -2928 33742 -2872
rect 33742 -2928 33762 -2872
rect 34678 -2868 34698 -2812
rect 34698 -2868 34722 -2812
rect 34722 -2868 34742 -2812
rect 34758 -2868 34778 -2812
rect 34778 -2868 34802 -2812
rect 34802 -2868 34822 -2812
rect 34678 -2872 34742 -2868
rect 34758 -2872 34822 -2868
rect 36878 -2812 36942 -2808
rect 36958 -2812 37022 -2808
rect 36878 -2868 36898 -2812
rect 36898 -2868 36922 -2812
rect 36922 -2868 36942 -2812
rect 36958 -2868 36978 -2812
rect 36978 -2868 37002 -2812
rect 37002 -2868 37022 -2812
rect 36878 -2872 36942 -2868
rect 36958 -2872 37022 -2868
rect 39078 -2812 39142 -2808
rect 39158 -2812 39222 -2808
rect 39078 -2868 39098 -2812
rect 39098 -2868 39122 -2812
rect 39122 -2868 39142 -2812
rect 39158 -2868 39178 -2812
rect 39178 -2868 39202 -2812
rect 39202 -2868 39222 -2812
rect 39078 -2872 39142 -2868
rect 39158 -2872 39222 -2868
rect 41278 -2812 41342 -2808
rect 41358 -2812 41422 -2808
rect 41278 -2868 41298 -2812
rect 41298 -2868 41322 -2812
rect 41322 -2868 41342 -2812
rect 41358 -2868 41378 -2812
rect 41378 -2868 41402 -2812
rect 41402 -2868 41422 -2812
rect 41278 -2872 41342 -2868
rect 41358 -2872 41422 -2868
rect 43478 -2812 43542 -2808
rect 43558 -2812 43622 -2808
rect 43478 -2868 43498 -2812
rect 43498 -2868 43522 -2812
rect 43522 -2868 43542 -2812
rect 43558 -2868 43578 -2812
rect 43578 -2868 43602 -2812
rect 43602 -2868 43622 -2812
rect 43478 -2872 43542 -2868
rect 43558 -2872 43622 -2868
rect 61838 -2872 61902 -2868
rect 61918 -2872 61982 -2868
rect 61998 -2872 62062 -2868
rect 33538 -2932 33602 -2928
rect 33618 -2932 33682 -2928
rect 33698 -2932 33762 -2928
rect 61838 -2928 61858 -2872
rect 61858 -2928 61882 -2872
rect 61882 -2928 61902 -2872
rect 61918 -2928 61938 -2872
rect 61938 -2928 61962 -2872
rect 61962 -2928 61982 -2872
rect 61998 -2928 62018 -2872
rect 62018 -2928 62042 -2872
rect 62042 -2928 62062 -2872
rect 61838 -2932 61902 -2928
rect 61918 -2932 61982 -2928
rect 61998 -2932 62062 -2928
rect -14092 -9212 -13708 -9208
rect -14092 -9988 -14088 -9212
rect -14088 -9988 -13712 -9212
rect -13712 -9988 -13708 -9212
rect -14092 -9992 -13708 -9988
rect 9638 -10272 9702 -10268
rect 9718 -10272 9782 -10268
rect 9798 -10272 9862 -10268
rect 9638 -10328 9658 -10272
rect 9658 -10328 9682 -10272
rect 9682 -10328 9702 -10272
rect 9718 -10328 9738 -10272
rect 9738 -10328 9762 -10272
rect 9762 -10328 9782 -10272
rect 9798 -10328 9818 -10272
rect 9818 -10328 9842 -10272
rect 9842 -10328 9862 -10272
rect 9638 -10332 9702 -10328
rect 9718 -10332 9782 -10328
rect 9798 -10332 9862 -10328
rect 35736 -10272 35800 -10268
rect 35816 -10272 35880 -10268
rect 35896 -10272 35960 -10268
rect 35736 -10328 35756 -10272
rect 35756 -10328 35780 -10272
rect 35780 -10328 35800 -10272
rect 35816 -10328 35836 -10272
rect 35836 -10328 35860 -10272
rect 35860 -10328 35880 -10272
rect 35896 -10328 35916 -10272
rect 35916 -10328 35940 -10272
rect 35940 -10328 35960 -10272
rect 35736 -10332 35800 -10328
rect 35816 -10332 35880 -10328
rect 35896 -10332 35960 -10328
rect 61838 -10272 61902 -10268
rect 61918 -10272 61982 -10268
rect 61998 -10272 62062 -10268
rect 61838 -10328 61858 -10272
rect 61858 -10328 61882 -10272
rect 61882 -10328 61902 -10272
rect 61918 -10328 61938 -10272
rect 61938 -10328 61962 -10272
rect 61962 -10328 61982 -10272
rect 61998 -10328 62018 -10272
rect 62018 -10328 62042 -10272
rect 62042 -10328 62062 -10272
rect 61838 -10332 61902 -10328
rect 61918 -10332 61982 -10328
rect 61998 -10332 62062 -10328
<< metal4 >>
rect -14220 11800 62300 12000
rect -14220 9722 -14020 11800
rect -14220 9658 -14152 9722
rect -14088 9658 -14020 9722
rect -14220 7400 -14020 9658
rect -10920 11252 -10780 11800
rect -10920 11188 -10882 11252
rect -10818 11188 -10780 11252
rect -10920 11172 -10780 11188
rect -10920 11108 -10882 11172
rect -10818 11108 -10780 11172
rect -10920 11092 -10780 11108
rect -10920 11028 -10882 11092
rect -10818 11028 -10780 11092
rect -10920 11012 -10780 11028
rect -10920 10948 -10882 11012
rect -10818 10948 -10780 11012
rect -10920 10932 -10780 10948
rect -10920 10868 -10882 10932
rect -10818 10868 -10780 10932
rect -10920 10852 -10780 10868
rect -10920 10788 -10882 10852
rect -10818 10788 -10780 10852
rect -10920 10772 -10780 10788
rect -10920 10708 -10882 10772
rect -10818 10708 -10780 10772
rect -10920 10692 -10780 10708
rect -10920 10628 -10882 10692
rect -10818 10628 -10780 10692
rect -10920 10612 -10780 10628
rect -10920 10548 -10882 10612
rect -10818 10548 -10780 10612
rect -8800 10581 -8600 11800
rect -10920 10532 -10780 10548
rect -10920 10468 -10882 10532
rect -10818 10468 -10780 10532
rect -10920 10452 -10780 10468
rect -10920 10388 -10882 10452
rect -10818 10388 -10780 10452
rect -10920 10372 -10780 10388
rect -10920 10308 -10882 10372
rect -10818 10308 -10780 10372
rect -10920 10292 -10780 10308
rect -10920 10228 -10882 10292
rect -10818 10228 -10780 10292
rect -10920 10212 -10780 10228
rect -10920 10148 -10882 10212
rect -10818 10148 -10780 10212
rect -8801 10542 -8600 10581
rect -8801 10478 -8772 10542
rect -8708 10478 -8600 10542
rect -8801 10462 -8600 10478
rect -8801 10398 -8772 10462
rect -8708 10398 -8600 10462
rect -8801 10382 -8600 10398
rect -8801 10318 -8772 10382
rect -8708 10318 -8600 10382
rect -8801 10302 -8600 10318
rect -8801 10238 -8772 10302
rect -8708 10238 -8600 10302
rect -8801 10199 -8600 10238
rect -10920 10132 -10780 10148
rect -10920 10068 -10882 10132
rect -10818 10068 -10780 10132
rect -10920 9722 -10780 10068
rect -10920 9658 -10882 9722
rect -10818 9658 -10780 9722
rect -10920 7580 -10780 9658
rect -8800 7500 -8600 10199
rect -3500 9272 -2800 9300
rect -3500 9128 -2972 9272
rect -2828 9128 -2800 9272
rect -3500 9100 -2800 9128
rect -7021 3240 -6899 3241
rect 4600 3240 4800 11800
rect -7021 3212 4800 3240
rect -7021 3148 -6992 3212
rect -6928 3148 4800 3212
rect -7021 3132 4800 3148
rect -7021 3068 -6992 3132
rect -6928 3068 4800 3132
rect -7021 3040 4800 3068
rect -7021 3039 -6899 3040
rect -2140 2540 -1400 2740
rect -1600 -2408 -1400 2540
rect 4600 400 4800 3040
rect 4600 352 5100 400
rect 4600 208 4698 352
rect 5002 208 5100 352
rect 4600 180 5100 208
rect -1600 -2472 -1532 -2408
rect -1468 -2472 -1400 -2408
rect -1600 -2488 -1400 -2472
rect -1600 -2552 -1532 -2488
rect -1468 -2552 -1400 -2488
rect -1600 -3180 -1400 -2552
rect 28039 -2800 28261 -2799
rect 30239 -2800 30461 -2799
rect 32439 -2800 32661 -2799
rect 34639 -2800 34861 -2799
rect 36839 -2800 37061 -2799
rect 39039 -2800 39261 -2799
rect 41239 -2800 41461 -2799
rect 43439 -2800 43661 -2799
rect 9300 -2808 62400 -2800
rect 9300 -2868 28078 -2808
rect 9300 -2932 9658 -2868
rect 9722 -2932 9738 -2868
rect 9802 -2932 9818 -2868
rect 9882 -2872 28078 -2868
rect 28142 -2872 28158 -2808
rect 28222 -2872 30278 -2808
rect 30342 -2872 30358 -2808
rect 30422 -2872 32478 -2808
rect 32542 -2872 32558 -2808
rect 32622 -2868 34678 -2808
rect 32622 -2872 33538 -2868
rect 9882 -2932 33538 -2872
rect 33602 -2932 33618 -2868
rect 33682 -2932 33698 -2868
rect 33762 -2872 34678 -2868
rect 34742 -2872 34758 -2808
rect 34822 -2872 36878 -2808
rect 36942 -2872 36958 -2808
rect 37022 -2872 39078 -2808
rect 39142 -2872 39158 -2808
rect 39222 -2872 41278 -2808
rect 41342 -2872 41358 -2808
rect 41422 -2872 43478 -2808
rect 43542 -2872 43558 -2808
rect 43622 -2868 62400 -2808
rect 43622 -2872 61838 -2868
rect 33762 -2932 61838 -2872
rect 61902 -2932 61918 -2868
rect 61982 -2932 61998 -2868
rect 62062 -2932 62400 -2868
rect 9300 -3000 62400 -2932
rect -14220 -3559 -14020 -3240
rect -2580 -3380 -1380 -3180
rect -1600 -3400 -1400 -3380
rect -14220 -3598 -13659 -3559
rect -14220 -3742 -14132 -3598
rect -13668 -3742 -13659 -3598
rect -14220 -3781 -13659 -3742
rect -14220 -9199 -14020 -3781
rect -14220 -9208 -13699 -9199
rect -14220 -9992 -14092 -9208
rect -13708 -9992 -13699 -9208
rect -14220 -10001 -13699 -9992
rect -14220 -10200 -14020 -10001
rect 9300 -10200 9600 -3000
rect 62200 -10200 62400 -3000
rect -14220 -10268 62400 -10200
rect -14220 -10332 9638 -10268
rect 9702 -10332 9718 -10268
rect 9782 -10332 9798 -10268
rect 9862 -10332 35736 -10268
rect 35800 -10332 35816 -10268
rect 35880 -10332 35896 -10268
rect 35960 -10332 61838 -10268
rect 61902 -10332 61918 -10268
rect 61982 -10332 61998 -10268
rect 62062 -10332 62400 -10268
rect -14220 -10400 62400 -10332
use XM_Rref  XM_Rref_0
timestamp 1663011646
transform 0 1 -13057 -1 0 -5305
box -1407 -1163 5019 21213
use XM_bjt  XM_bjt_0
timestamp 1663011646
transform 1 0 -2070 0 1 -2620
box 0 0 6492 9068
use XM_bjt_out  XM_bjt_out_0
timestamp 1663011646
transform 1 0 -2070 0 1 6780
box 0 0 6492 3916
use XM_current_gate_with_dummy  XM_current_gate_with_dummy_0
timestamp 1663011646
transform 1 0 4524 0 1 -1712
box 0 -924 4660 1954
use XM_feedbackmir2  XM_feedbackmir2_0
timestamp 1663011646
transform 1 0 -10768 0 1 9846
box -140 -160 2080 1600
use XM_feedbackmir  XM_feedbackmir_0
timestamp 1663011646
transform 1 0 -13500 0 1 8386
box -700 -500 2900 3100
use XM_otabias_nmos  XM_otabias_nmos_0
timestamp 1663011646
transform 1 0 -7877 0 1 9671
box -43 -43 1129 1295
use XM_otabias_pmos  XM_otabias_pmos_0
timestamp 1663011646
transform 1 0 -10817 0 1 8939
box -53 -53 1571 879
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1663011646
transform 1 0 26905 0 1 -3003
box -17526 -7326 35426 14926
use XM_pdn  XM_pdn_0
timestamp 1663011646
transform 1 0 -8785 0 1 9133
box -53 -708 5500 1206
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1663011646
transform 1 0 -8840 0 1 1874
box -5380 594 6766 6403
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_1
timestamp 1663011646
transform 1 0 -8840 0 1 -4044
box -5380 594 6766 6403
use sky130_fd_pr__res_high_po_1p41_6ZUZ5C  sky130_fd_pr__res_high_po_1p41_6ZUZ5C_0
timestamp 1663011646
transform 1 0 -8623 0 1 7103
box -297 -1398 297 1398
use sky130_fd_pr__res_high_po_1p41_GWJZ59  sky130_fd_pr__res_high_po_1p41_GWJZ59_0
timestamp 1663011646
transform 0 1 -3232 -1 0 -3669
box -297 -10988 297 10988
use sky130_fd_pr__res_high_po_1p41_HX7ZEK  sky130_fd_pr__res_high_po_1p41_HX7ZEK_0
timestamp 1663011646
transform 0 1 3187 -1 0 -3015
box -297 -5338 297 5338
use sky130_fd_pr__res_high_po_1p41_S8KB58  sky130_fd_pr__res_high_po_1p41_S8KB58_0
timestamp 1663011646
transform 0 1 -3253 -1 0 11177
box -297 -4827 297 4827
<< labels >>
flabel metal2 s -9540 5700 -9480 7680 0 FreeSans 1000 0 0 0 vb
port 1 nsew
flabel metal3 s -8760 8740 -8200 8840 0 FreeSans 1000 0 0 0 vgate
port 2 nsew
flabel metal2 s 1160 8800 1380 11100 0 FreeSans 1000 0 0 0 vbe3
port 3 nsew
flabel metal1 s -9200 -2991 -9100 5271 0 FreeSans 1000 0 0 0 Vota_bias1
port 4 nsew
flabel metal3 s 6920 -3800 7040 -1540 0 FreeSans 2000 0 0 0 vd4
port 5 nsew
flabel metal2 s 6420 320 6600 4600 0 FreeSans 4000 0 0 0 voutb2
port 6 nsew
flabel metal1 s -8700 8200 -4700 8400 0 FreeSans 4000 0 0 0 vbneg
port 7 nsew
flabel metal3 s 30200 4260 30500 12600 0 FreeSans 4000 0 0 0 Iout0
port 8 nsew
flabel metal4 s -14220 9760 -14020 12000 0 FreeSans 4000 0 0 0 VDD
port 9 nsew
flabel metal4 s -14220 -9200 -14020 -3780 0 FreeSans 4000 0 0 0 VSS
port 10 nsew
flabel metal3 s 32400 4260 32700 12600 0 FreeSans 4000 0 0 0 Iout1
port 11 nsew
flabel metal3 s 34600 4260 34900 12600 0 FreeSans 4000 0 0 0 Iout2
port 12 nsew
flabel metal3 s -8500 10860 -8380 12540 0 FreeSans 4000 0 0 0 porst
port 13 nsew
flabel metal2 s -7900 11120 -7700 12500 0 FreeSans 2000 0 0 0 vbg
port 14 nsew
flabel metal3 s 36800 4260 37100 12600 0 FreeSans 4000 0 0 0 Iout3
port 15 nsew
flabel metal3 s 39000 4260 39300 12600 0 FreeSans 4000 0 0 0 Iout4
port 16 nsew
flabel metal3 s 41200 4260 41500 12600 0 FreeSans 4000 0 0 0 Iout5
port 17 nsew
flabel metal3 s 43400 4260 43700 12600 0 FreeSans 4000 0 0 0 Iout6
port 18 nsew
<< end >>
