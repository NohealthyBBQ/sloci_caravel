magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -586 -669 586 669
<< nmoslvt >>
rect -400 -469 400 531
<< ndiff >>
rect -458 490 -400 531
rect -458 456 -446 490
rect -412 456 -400 490
rect -458 422 -400 456
rect -458 388 -446 422
rect -412 388 -400 422
rect -458 354 -400 388
rect -458 320 -446 354
rect -412 320 -400 354
rect -458 286 -400 320
rect -458 252 -446 286
rect -412 252 -400 286
rect -458 218 -400 252
rect -458 184 -446 218
rect -412 184 -400 218
rect -458 150 -400 184
rect -458 116 -446 150
rect -412 116 -400 150
rect -458 82 -400 116
rect -458 48 -446 82
rect -412 48 -400 82
rect -458 14 -400 48
rect -458 -20 -446 14
rect -412 -20 -400 14
rect -458 -54 -400 -20
rect -458 -88 -446 -54
rect -412 -88 -400 -54
rect -458 -122 -400 -88
rect -458 -156 -446 -122
rect -412 -156 -400 -122
rect -458 -190 -400 -156
rect -458 -224 -446 -190
rect -412 -224 -400 -190
rect -458 -258 -400 -224
rect -458 -292 -446 -258
rect -412 -292 -400 -258
rect -458 -326 -400 -292
rect -458 -360 -446 -326
rect -412 -360 -400 -326
rect -458 -394 -400 -360
rect -458 -428 -446 -394
rect -412 -428 -400 -394
rect -458 -469 -400 -428
rect 400 490 458 531
rect 400 456 412 490
rect 446 456 458 490
rect 400 422 458 456
rect 400 388 412 422
rect 446 388 458 422
rect 400 354 458 388
rect 400 320 412 354
rect 446 320 458 354
rect 400 286 458 320
rect 400 252 412 286
rect 446 252 458 286
rect 400 218 458 252
rect 400 184 412 218
rect 446 184 458 218
rect 400 150 458 184
rect 400 116 412 150
rect 446 116 458 150
rect 400 82 458 116
rect 400 48 412 82
rect 446 48 458 82
rect 400 14 458 48
rect 400 -20 412 14
rect 446 -20 458 14
rect 400 -54 458 -20
rect 400 -88 412 -54
rect 446 -88 458 -54
rect 400 -122 458 -88
rect 400 -156 412 -122
rect 446 -156 458 -122
rect 400 -190 458 -156
rect 400 -224 412 -190
rect 446 -224 458 -190
rect 400 -258 458 -224
rect 400 -292 412 -258
rect 446 -292 458 -258
rect 400 -326 458 -292
rect 400 -360 412 -326
rect 446 -360 458 -326
rect 400 -394 458 -360
rect 400 -428 412 -394
rect 446 -428 458 -394
rect 400 -469 458 -428
<< ndiffc >>
rect -446 456 -412 490
rect -446 388 -412 422
rect -446 320 -412 354
rect -446 252 -412 286
rect -446 184 -412 218
rect -446 116 -412 150
rect -446 48 -412 82
rect -446 -20 -412 14
rect -446 -88 -412 -54
rect -446 -156 -412 -122
rect -446 -224 -412 -190
rect -446 -292 -412 -258
rect -446 -360 -412 -326
rect -446 -428 -412 -394
rect 412 456 446 490
rect 412 388 446 422
rect 412 320 446 354
rect 412 252 446 286
rect 412 184 446 218
rect 412 116 446 150
rect 412 48 446 82
rect 412 -20 446 14
rect 412 -88 446 -54
rect 412 -156 446 -122
rect 412 -224 446 -190
rect 412 -292 446 -258
rect 412 -360 446 -326
rect 412 -428 446 -394
<< psubdiff >>
rect -560 609 560 643
rect -560 -609 -526 609
rect 526 -609 560 609
rect -560 -643 560 -609
<< poly >>
rect -400 531 400 557
rect -400 -507 400 -469
rect -400 -541 -357 -507
rect -323 -541 -289 -507
rect -255 -541 -221 -507
rect -187 -541 -153 -507
rect -119 -541 -85 -507
rect -51 -541 -17 -507
rect 17 -541 51 -507
rect 85 -541 119 -507
rect 153 -541 187 -507
rect 221 -541 255 -507
rect 289 -541 323 -507
rect 357 -541 400 -507
rect -400 -557 400 -541
<< polycont >>
rect -357 -541 -323 -507
rect -289 -541 -255 -507
rect -221 -541 -187 -507
rect -153 -541 -119 -507
rect -85 -541 -51 -507
rect -17 -541 17 -507
rect 51 -541 85 -507
rect 119 -541 153 -507
rect 187 -541 221 -507
rect 255 -541 289 -507
rect 323 -541 357 -507
<< locali >>
rect -560 609 560 643
rect -560 -609 -526 609
rect -446 516 -412 535
rect -446 444 -412 456
rect -446 372 -412 388
rect -446 300 -412 320
rect -446 228 -412 252
rect -446 156 -412 184
rect -446 84 -412 116
rect -446 14 -412 48
rect -446 -54 -412 -22
rect -446 -122 -412 -94
rect -446 -190 -412 -166
rect -446 -258 -412 -238
rect -446 -326 -412 -310
rect -446 -394 -412 -382
rect -446 -473 -412 -454
rect 412 516 446 535
rect 412 444 446 456
rect 412 372 446 388
rect 412 300 446 320
rect 412 228 446 252
rect 412 156 446 184
rect 412 84 446 116
rect 412 14 446 48
rect 412 -54 446 -22
rect 412 -122 446 -94
rect 412 -190 446 -166
rect 412 -258 446 -238
rect 412 -326 446 -310
rect 412 -394 446 -382
rect 412 -473 446 -454
rect -400 -541 -377 -507
rect -323 -541 -305 -507
rect -255 -541 -233 -507
rect -187 -541 -161 -507
rect -119 -541 -89 -507
rect -51 -541 -17 -507
rect 17 -541 51 -507
rect 89 -541 119 -507
rect 161 -541 187 -507
rect 233 -541 255 -507
rect 305 -541 323 -507
rect 377 -541 400 -507
rect 526 -609 560 609
rect -560 -643 560 -609
<< viali >>
rect -446 490 -412 516
rect -446 482 -412 490
rect -446 422 -412 444
rect -446 410 -412 422
rect -446 354 -412 372
rect -446 338 -412 354
rect -446 286 -412 300
rect -446 266 -412 286
rect -446 218 -412 228
rect -446 194 -412 218
rect -446 150 -412 156
rect -446 122 -412 150
rect -446 82 -412 84
rect -446 50 -412 82
rect -446 -20 -412 12
rect -446 -22 -412 -20
rect -446 -88 -412 -60
rect -446 -94 -412 -88
rect -446 -156 -412 -132
rect -446 -166 -412 -156
rect -446 -224 -412 -204
rect -446 -238 -412 -224
rect -446 -292 -412 -276
rect -446 -310 -412 -292
rect -446 -360 -412 -348
rect -446 -382 -412 -360
rect -446 -428 -412 -420
rect -446 -454 -412 -428
rect 412 490 446 516
rect 412 482 446 490
rect 412 422 446 444
rect 412 410 446 422
rect 412 354 446 372
rect 412 338 446 354
rect 412 286 446 300
rect 412 266 446 286
rect 412 218 446 228
rect 412 194 446 218
rect 412 150 446 156
rect 412 122 446 150
rect 412 82 446 84
rect 412 50 446 82
rect 412 -20 446 12
rect 412 -22 446 -20
rect 412 -88 446 -60
rect 412 -94 446 -88
rect 412 -156 446 -132
rect 412 -166 446 -156
rect 412 -224 446 -204
rect 412 -238 446 -224
rect 412 -292 446 -276
rect 412 -310 446 -292
rect 412 -360 446 -348
rect 412 -382 446 -360
rect 412 -428 446 -420
rect 412 -454 446 -428
rect -377 -541 -357 -507
rect -357 -541 -343 -507
rect -305 -541 -289 -507
rect -289 -541 -271 -507
rect -233 -541 -221 -507
rect -221 -541 -199 -507
rect -161 -541 -153 -507
rect -153 -541 -127 -507
rect -89 -541 -85 -507
rect -85 -541 -55 -507
rect -17 -541 17 -507
rect 55 -541 85 -507
rect 85 -541 89 -507
rect 127 -541 153 -507
rect 153 -541 161 -507
rect 199 -541 221 -507
rect 221 -541 233 -507
rect 271 -541 289 -507
rect 289 -541 305 -507
rect 343 -541 357 -507
rect 357 -541 377 -507
<< metal1 >>
rect -452 516 -406 531
rect -452 482 -446 516
rect -412 482 -406 516
rect -452 444 -406 482
rect -452 410 -446 444
rect -412 410 -406 444
rect -452 372 -406 410
rect -452 338 -446 372
rect -412 338 -406 372
rect -452 300 -406 338
rect -452 266 -446 300
rect -412 266 -406 300
rect -452 228 -406 266
rect -452 194 -446 228
rect -412 194 -406 228
rect -452 156 -406 194
rect -452 122 -446 156
rect -412 122 -406 156
rect -452 84 -406 122
rect -452 50 -446 84
rect -412 50 -406 84
rect -452 12 -406 50
rect -452 -22 -446 12
rect -412 -22 -406 12
rect -452 -60 -406 -22
rect -452 -94 -446 -60
rect -412 -94 -406 -60
rect -452 -132 -406 -94
rect -452 -166 -446 -132
rect -412 -166 -406 -132
rect -452 -204 -406 -166
rect -452 -238 -446 -204
rect -412 -238 -406 -204
rect -452 -276 -406 -238
rect -452 -310 -446 -276
rect -412 -310 -406 -276
rect -452 -348 -406 -310
rect -452 -382 -446 -348
rect -412 -382 -406 -348
rect -452 -420 -406 -382
rect -452 -454 -446 -420
rect -412 -454 -406 -420
rect -452 -469 -406 -454
rect 406 516 452 531
rect 406 482 412 516
rect 446 482 452 516
rect 406 444 452 482
rect 406 410 412 444
rect 446 410 452 444
rect 406 372 452 410
rect 406 338 412 372
rect 446 338 452 372
rect 406 300 452 338
rect 406 266 412 300
rect 446 266 452 300
rect 406 228 452 266
rect 406 194 412 228
rect 446 194 452 228
rect 406 156 452 194
rect 406 122 412 156
rect 446 122 452 156
rect 406 84 452 122
rect 406 50 412 84
rect 446 50 452 84
rect 406 12 452 50
rect 406 -22 412 12
rect 446 -22 452 12
rect 406 -60 452 -22
rect 406 -94 412 -60
rect 446 -94 452 -60
rect 406 -132 452 -94
rect 406 -166 412 -132
rect 446 -166 452 -132
rect 406 -204 452 -166
rect 406 -238 412 -204
rect 446 -238 452 -204
rect 406 -276 452 -238
rect 406 -310 412 -276
rect 446 -310 452 -276
rect 406 -348 452 -310
rect 406 -382 412 -348
rect 446 -382 452 -348
rect 406 -420 452 -382
rect 406 -454 412 -420
rect 446 -454 452 -420
rect 406 -469 452 -454
rect -396 -507 396 -501
rect -396 -541 -377 -507
rect -343 -541 -305 -507
rect -271 -541 -233 -507
rect -199 -541 -161 -507
rect -127 -541 -89 -507
rect -55 -541 -17 -507
rect 17 -541 55 -507
rect 89 -541 127 -507
rect 161 -541 199 -507
rect 233 -541 271 -507
rect 305 -541 343 -507
rect 377 -541 396 -507
rect -396 -547 396 -541
<< properties >>
string FIXED_BBOX -543 -626 543 626
<< end >>
