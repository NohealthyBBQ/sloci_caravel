magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 33895 33129 34005 33155
rect 33895 33095 33933 33129
rect 33967 33095 34005 33129
rect 33895 33070 34005 33095
rect 55194 32310 55348 32350
rect 33260 32123 33380 32155
rect 33260 32089 33303 32123
rect 33337 32089 33380 32123
rect 33260 32051 33380 32089
rect 33260 32017 33303 32051
rect 33337 32017 33380 32051
rect 33260 31990 33380 32017
rect 52140 31536 52255 31580
rect 52140 31502 52178 31536
rect 52212 31502 52255 31536
rect 52140 31464 52255 31502
rect 52140 31430 52178 31464
rect 52212 31430 52255 31464
rect 52140 31392 52255 31430
rect 52140 31358 52178 31392
rect 52212 31358 52255 31392
rect 52140 31320 52255 31358
rect 52140 31286 52178 31320
rect 52212 31286 52255 31320
rect 52140 31248 52255 31286
rect 36440 31187 36900 31220
rect 36440 31153 36473 31187
rect 36507 31153 36545 31187
rect 36579 31153 36617 31187
rect 36651 31153 36689 31187
rect 36723 31153 36761 31187
rect 36795 31153 36833 31187
rect 36867 31153 36900 31187
rect 52140 31214 52178 31248
rect 52212 31214 52255 31248
rect 52140 31175 52255 31214
rect 36440 31120 36900 31153
rect 55184 29702 55338 29742
rect 55174 27882 55328 27922
rect 52135 26413 52250 26455
rect 52135 26379 52173 26413
rect 52207 26379 52250 26413
rect 52135 26341 52250 26379
rect 52135 26307 52173 26341
rect 52207 26307 52250 26341
rect 52135 26269 52250 26307
rect 52135 26235 52173 26269
rect 52207 26235 52250 26269
rect 52135 26197 52250 26235
rect 52135 26163 52173 26197
rect 52207 26163 52250 26197
rect 52135 26125 52250 26163
rect 52135 26091 52173 26125
rect 52207 26091 52250 26125
rect 52135 26050 52250 26091
rect 34160 25810 36370 25850
rect 36420 25580 36940 25590
rect 33670 25567 36940 25580
rect 33670 25540 36447 25567
rect 36420 25533 36447 25540
rect 36481 25533 36519 25567
rect 36553 25533 36591 25567
rect 36625 25533 36663 25567
rect 36697 25533 36735 25567
rect 36769 25533 36807 25567
rect 36841 25533 36879 25567
rect 36913 25533 36940 25567
rect 36420 25510 36940 25533
rect 55178 25280 55332 25320
rect 32925 24439 33320 24480
rect 32925 24405 32959 24439
rect 32993 24405 33031 24439
rect 33065 24405 33103 24439
rect 33137 24405 33175 24439
rect 33209 24405 33247 24439
rect 33281 24405 33320 24439
rect 32925 24370 33320 24405
<< viali >>
rect 33933 33095 33967 33129
rect 33303 32089 33337 32123
rect 33303 32017 33337 32051
rect 52178 31502 52212 31536
rect 52178 31430 52212 31464
rect 52178 31358 52212 31392
rect 52178 31286 52212 31320
rect 36473 31153 36507 31187
rect 36545 31153 36579 31187
rect 36617 31153 36651 31187
rect 36689 31153 36723 31187
rect 36761 31153 36795 31187
rect 36833 31153 36867 31187
rect 52178 31214 52212 31248
rect 52173 26379 52207 26413
rect 52173 26307 52207 26341
rect 52173 26235 52207 26269
rect 52173 26163 52207 26197
rect 52173 26091 52207 26125
rect 36447 25533 36481 25567
rect 36519 25533 36553 25567
rect 36591 25533 36625 25567
rect 36663 25533 36697 25567
rect 36735 25533 36769 25567
rect 36807 25533 36841 25567
rect 36879 25533 36913 25567
rect 32959 24405 32993 24439
rect 33031 24405 33065 24439
rect 33103 24405 33137 24439
rect 33175 24405 33209 24439
rect 33247 24405 33281 24439
<< metal1 >>
rect 46750 37650 46800 38020
rect 46210 37580 46800 37650
rect 33895 33138 34005 33155
rect 33895 33086 33924 33138
rect 33976 33086 34005 33138
rect 33895 33070 34005 33086
rect 33475 32875 33520 33000
rect 33590 32988 33665 33000
rect 33590 32936 33601 32988
rect 33653 32936 33665 32988
rect 33590 32925 33665 32936
rect 33455 32863 33530 32875
rect 33455 32811 33466 32863
rect 33518 32811 33530 32863
rect 33455 32800 33530 32811
rect 33605 32800 33650 32925
rect 33730 32875 33775 33000
rect 33845 32988 33920 33000
rect 33845 32936 33856 32988
rect 33908 32936 33920 32988
rect 33845 32925 33920 32936
rect 33715 32863 33790 32875
rect 33715 32811 33726 32863
rect 33778 32811 33790 32863
rect 33715 32800 33790 32811
rect 33860 32800 33905 32925
rect 33520 32743 33865 32755
rect 33520 32715 33796 32743
rect 33780 32691 33796 32715
rect 33848 32691 33865 32743
rect 33780 32210 33865 32691
rect 36090 32690 36320 32760
rect 46210 32690 46280 37580
rect 47720 36710 47775 37940
rect 48190 36710 48240 38290
rect 47700 36695 47790 36710
rect 47700 36643 47719 36695
rect 47771 36643 47790 36695
rect 47700 36631 47790 36643
rect 47700 36579 47719 36631
rect 47771 36579 47790 36631
rect 47700 36567 47790 36579
rect 47700 36515 47719 36567
rect 47771 36515 47790 36567
rect 47700 36500 47790 36515
rect 48170 36695 48260 36710
rect 48170 36643 48189 36695
rect 48241 36643 48260 36695
rect 48170 36631 48260 36643
rect 48170 36579 48189 36631
rect 48241 36579 48260 36631
rect 48170 36567 48260 36579
rect 48170 36515 48189 36567
rect 48241 36515 48260 36567
rect 48170 36500 48260 36515
rect 33260 32128 33380 32155
rect 33260 32076 33294 32128
rect 33346 32076 33380 32128
rect 33260 32064 33380 32076
rect 33260 32012 33294 32064
rect 33346 32012 33380 32064
rect 33260 31990 33380 32012
rect 35740 30959 35980 31000
rect 35740 30651 35770 30959
rect 35950 30651 35980 30959
rect 35740 30640 35980 30651
rect 35580 30580 35980 30640
rect 35761 27556 35862 27557
rect 35620 27495 35862 27556
rect 35761 27001 35862 27495
rect 35761 26949 35785 27001
rect 35837 26949 35862 27001
rect 35761 26937 35862 26949
rect 35761 26885 35785 26937
rect 35837 26885 35862 26937
rect 35761 26873 35862 26885
rect 35761 26821 35785 26873
rect 35837 26821 35862 26873
rect 35761 26809 35862 26821
rect 35761 26757 35785 26809
rect 35837 26757 35862 26809
rect 35761 26745 35862 26757
rect 35761 26693 35785 26745
rect 35837 26693 35862 26745
rect 35761 26681 35862 26693
rect 35761 26629 35785 26681
rect 35837 26629 35862 26681
rect 35761 26603 35862 26629
rect 36090 25345 36160 32690
rect 36440 31187 36900 31220
rect 36440 31153 36473 31187
rect 36507 31176 36545 31187
rect 36579 31176 36617 31187
rect 36651 31176 36689 31187
rect 36723 31176 36761 31187
rect 36795 31176 36833 31187
rect 36536 31153 36545 31176
rect 36440 31124 36484 31153
rect 36536 31124 36548 31153
rect 36600 31124 36612 31176
rect 36664 31124 36676 31176
rect 36728 31124 36740 31176
rect 36795 31153 36804 31176
rect 36867 31153 36900 31187
rect 46335 31170 46440 31580
rect 36792 31124 36804 31153
rect 36856 31124 36900 31153
rect 36440 31100 36900 31124
rect 50680 31080 50730 37490
rect 57390 36205 57750 36265
rect 59485 36205 59860 36265
rect 61580 36205 61955 36265
rect 63670 36205 64910 36265
rect 57365 35845 57745 35905
rect 59490 35845 59865 35905
rect 61585 35845 61960 35905
rect 63690 35845 64655 35905
rect 57355 35305 57730 35365
rect 59465 35305 59840 35365
rect 61595 35305 61970 35365
rect 63660 35305 64405 35365
rect 57380 34715 57755 34775
rect 59460 34715 59835 34775
rect 61570 34715 61945 34775
rect 63655 34715 64140 34775
rect 57385 33805 57760 33865
rect 59460 33805 59835 33865
rect 61555 33805 61930 33865
rect 63700 33805 63905 33865
rect 52140 31536 52255 31580
rect 52140 31529 52178 31536
rect 52212 31529 52255 31536
rect 52140 31477 52169 31529
rect 52221 31477 52255 31529
rect 52140 31465 52255 31477
rect 52140 31413 52169 31465
rect 52221 31413 52255 31465
rect 52140 31401 52255 31413
rect 52140 31349 52169 31401
rect 52221 31349 52255 31401
rect 52140 31337 52255 31349
rect 52140 31285 52169 31337
rect 52221 31285 52255 31337
rect 52140 31273 52255 31285
rect 52140 31221 52169 31273
rect 52221 31221 52255 31273
rect 52140 31214 52178 31221
rect 52212 31214 52255 31221
rect 52140 31175 52255 31214
rect 55108 31074 56370 31134
rect 56292 31042 56370 31074
rect 56290 26556 56366 26586
rect 55094 26496 56366 26556
rect 52135 26438 52250 26455
rect 52135 26386 52164 26438
rect 52216 26386 52250 26438
rect 52135 26379 52173 26386
rect 52207 26379 52250 26386
rect 52135 26374 52250 26379
rect 52135 26322 52164 26374
rect 52216 26322 52250 26374
rect 52135 26310 52173 26322
rect 52207 26310 52250 26322
rect 52135 26258 52164 26310
rect 52216 26258 52250 26310
rect 52135 26246 52173 26258
rect 52207 26246 52250 26258
rect 52135 26194 52164 26246
rect 52216 26194 52250 26246
rect 52135 26182 52173 26194
rect 52207 26182 52250 26194
rect 52135 26130 52164 26182
rect 52216 26130 52250 26182
rect 52135 26125 52250 26130
rect 52135 26118 52173 26125
rect 52207 26118 52250 26125
rect 52135 26066 52164 26118
rect 52216 26066 52250 26118
rect 52135 26050 52250 26066
rect 36420 25567 36940 25590
rect 36420 25536 36447 25567
rect 36481 25536 36519 25567
rect 36553 25536 36591 25567
rect 36625 25536 36663 25567
rect 36697 25536 36735 25567
rect 36769 25536 36807 25567
rect 36841 25536 36879 25567
rect 36913 25536 36940 25567
rect 36420 25484 36430 25536
rect 36482 25484 36494 25536
rect 36553 25533 36558 25536
rect 36802 25533 36807 25536
rect 36546 25484 36558 25533
rect 36610 25484 36622 25533
rect 36674 25484 36686 25533
rect 36738 25484 36750 25533
rect 36802 25484 36814 25533
rect 36866 25484 36878 25536
rect 36930 25484 36940 25536
rect 36420 25470 36940 25484
rect 36045 25304 36160 25345
rect 36045 25252 36074 25304
rect 36126 25252 36160 25304
rect 36045 25240 36160 25252
rect 36045 25188 36074 25240
rect 36126 25188 36160 25240
rect 36045 25176 36160 25188
rect 36045 25124 36074 25176
rect 36126 25124 36160 25176
rect 36045 25112 36160 25124
rect 36045 25060 36074 25112
rect 36126 25060 36160 25112
rect 36045 25020 36160 25060
rect 32925 24448 33320 24480
rect 32925 24439 32966 24448
rect 32925 24405 32959 24439
rect 32925 24396 32966 24405
rect 33018 24396 33030 24448
rect 33082 24396 33094 24448
rect 33146 24396 33158 24448
rect 33210 24396 33222 24448
rect 33274 24439 33320 24448
rect 33281 24405 33320 24439
rect 33274 24396 33320 24405
rect 32925 24370 33320 24396
rect 36090 24050 36160 25020
rect 36090 23980 36400 24050
rect 63845 23825 63905 33805
rect 57370 23765 57745 23825
rect 59445 23765 59820 23825
rect 61580 23765 61955 23825
rect 63585 23765 63905 23825
rect 64080 22915 64140 34715
rect 57350 22855 57725 22915
rect 59460 22855 59835 22915
rect 61575 22855 61950 22915
rect 63635 22855 64140 22915
rect 64345 22325 64405 35305
rect 57370 22265 57745 22325
rect 59460 22265 59835 22325
rect 61575 22265 61950 22325
rect 63645 22265 64405 22325
rect 64595 21785 64655 35845
rect 57370 21725 57745 21785
rect 59475 21725 59850 21785
rect 61565 21725 61940 21785
rect 63700 21725 64655 21785
rect 64850 21425 64910 36205
rect 57360 21365 57735 21425
rect 59480 21365 59855 21425
rect 61570 21365 61945 21425
rect 63690 21365 64910 21425
<< via1 >>
rect 33924 33129 33976 33138
rect 33924 33095 33933 33129
rect 33933 33095 33967 33129
rect 33967 33095 33976 33129
rect 33924 33086 33976 33095
rect 33601 32936 33653 32988
rect 33466 32811 33518 32863
rect 33856 32936 33908 32988
rect 33726 32811 33778 32863
rect 33796 32691 33848 32743
rect 47719 36643 47771 36695
rect 47719 36579 47771 36631
rect 47719 36515 47771 36567
rect 48189 36643 48241 36695
rect 48189 36579 48241 36631
rect 48189 36515 48241 36567
rect 33294 32123 33346 32128
rect 33294 32089 33303 32123
rect 33303 32089 33337 32123
rect 33337 32089 33346 32123
rect 33294 32076 33346 32089
rect 33294 32051 33346 32064
rect 33294 32017 33303 32051
rect 33303 32017 33337 32051
rect 33337 32017 33346 32051
rect 33294 32012 33346 32017
rect 35770 30651 35950 30959
rect 35785 26949 35837 27001
rect 35785 26885 35837 26937
rect 35785 26821 35837 26873
rect 35785 26757 35837 26809
rect 35785 26693 35837 26745
rect 35785 26629 35837 26681
rect 36484 31153 36507 31176
rect 36507 31153 36536 31176
rect 36548 31153 36579 31176
rect 36579 31153 36600 31176
rect 36484 31124 36536 31153
rect 36548 31124 36600 31153
rect 36612 31153 36617 31176
rect 36617 31153 36651 31176
rect 36651 31153 36664 31176
rect 36612 31124 36664 31153
rect 36676 31153 36689 31176
rect 36689 31153 36723 31176
rect 36723 31153 36728 31176
rect 36676 31124 36728 31153
rect 36740 31153 36761 31176
rect 36761 31153 36792 31176
rect 36804 31153 36833 31176
rect 36833 31153 36856 31176
rect 36740 31124 36792 31153
rect 36804 31124 36856 31153
rect 52169 31502 52178 31529
rect 52178 31502 52212 31529
rect 52212 31502 52221 31529
rect 52169 31477 52221 31502
rect 52169 31464 52221 31465
rect 52169 31430 52178 31464
rect 52178 31430 52212 31464
rect 52212 31430 52221 31464
rect 52169 31413 52221 31430
rect 52169 31392 52221 31401
rect 52169 31358 52178 31392
rect 52178 31358 52212 31392
rect 52212 31358 52221 31392
rect 52169 31349 52221 31358
rect 52169 31320 52221 31337
rect 52169 31286 52178 31320
rect 52178 31286 52212 31320
rect 52212 31286 52221 31320
rect 52169 31285 52221 31286
rect 52169 31248 52221 31273
rect 52169 31221 52178 31248
rect 52178 31221 52212 31248
rect 52212 31221 52221 31248
rect 52164 26413 52216 26438
rect 52164 26386 52173 26413
rect 52173 26386 52207 26413
rect 52207 26386 52216 26413
rect 52164 26341 52216 26374
rect 52164 26322 52173 26341
rect 52173 26322 52207 26341
rect 52207 26322 52216 26341
rect 52164 26307 52173 26310
rect 52173 26307 52207 26310
rect 52207 26307 52216 26310
rect 52164 26269 52216 26307
rect 52164 26258 52173 26269
rect 52173 26258 52207 26269
rect 52207 26258 52216 26269
rect 52164 26235 52173 26246
rect 52173 26235 52207 26246
rect 52207 26235 52216 26246
rect 52164 26197 52216 26235
rect 52164 26194 52173 26197
rect 52173 26194 52207 26197
rect 52207 26194 52216 26197
rect 52164 26163 52173 26182
rect 52173 26163 52207 26182
rect 52207 26163 52216 26182
rect 52164 26130 52216 26163
rect 52164 26091 52173 26118
rect 52173 26091 52207 26118
rect 52207 26091 52216 26118
rect 52164 26066 52216 26091
rect 36430 25533 36447 25536
rect 36447 25533 36481 25536
rect 36481 25533 36482 25536
rect 36430 25484 36482 25533
rect 36494 25533 36519 25536
rect 36519 25533 36546 25536
rect 36558 25533 36591 25536
rect 36591 25533 36610 25536
rect 36622 25533 36625 25536
rect 36625 25533 36663 25536
rect 36663 25533 36674 25536
rect 36686 25533 36697 25536
rect 36697 25533 36735 25536
rect 36735 25533 36738 25536
rect 36750 25533 36769 25536
rect 36769 25533 36802 25536
rect 36814 25533 36841 25536
rect 36841 25533 36866 25536
rect 36494 25484 36546 25533
rect 36558 25484 36610 25533
rect 36622 25484 36674 25533
rect 36686 25484 36738 25533
rect 36750 25484 36802 25533
rect 36814 25484 36866 25533
rect 36878 25533 36879 25536
rect 36879 25533 36913 25536
rect 36913 25533 36930 25536
rect 36878 25484 36930 25533
rect 36074 25252 36126 25304
rect 36074 25188 36126 25240
rect 36074 25124 36126 25176
rect 36074 25060 36126 25112
rect 32966 24439 33018 24448
rect 32966 24405 32993 24439
rect 32993 24405 33018 24439
rect 32966 24396 33018 24405
rect 33030 24439 33082 24448
rect 33030 24405 33031 24439
rect 33031 24405 33065 24439
rect 33065 24405 33082 24439
rect 33030 24396 33082 24405
rect 33094 24439 33146 24448
rect 33094 24405 33103 24439
rect 33103 24405 33137 24439
rect 33137 24405 33146 24439
rect 33094 24396 33146 24405
rect 33158 24439 33210 24448
rect 33158 24405 33175 24439
rect 33175 24405 33209 24439
rect 33209 24405 33210 24439
rect 33158 24396 33210 24405
rect 33222 24439 33274 24448
rect 33222 24405 33247 24439
rect 33247 24405 33274 24439
rect 33222 24396 33274 24405
<< metal2 >>
rect 43710 38248 44220 38270
rect 43710 37952 43737 38248
rect 44193 37952 44220 38248
rect 43710 37930 44220 37952
rect 54790 37158 63380 37200
rect 54790 36800 54812 37158
rect 47700 36695 47790 36710
rect 47700 36673 47719 36695
rect 47771 36673 47790 36695
rect 47700 36617 47717 36673
rect 47773 36617 47790 36673
rect 47700 36593 47719 36617
rect 47771 36593 47790 36617
rect 47700 36537 47717 36593
rect 47773 36537 47790 36593
rect 47700 36515 47719 36537
rect 47771 36515 47790 36537
rect 47700 36500 47790 36515
rect 48170 36695 48260 36710
rect 48170 36673 48189 36695
rect 48241 36673 48260 36695
rect 48170 36617 48187 36673
rect 48243 36617 48260 36673
rect 48170 36593 48189 36617
rect 48241 36593 48260 36617
rect 54785 36622 54812 36800
rect 55188 36622 63380 37158
rect 54785 36600 63380 36622
rect 48170 36537 48187 36593
rect 48243 36537 48260 36593
rect 48170 36515 48189 36537
rect 48241 36515 48260 36537
rect 48170 36500 48260 36515
rect 55046 36460 55170 36462
rect 34240 36430 45110 36460
rect 34240 36428 45430 36430
rect 34240 36052 34279 36428
rect 34495 36393 45430 36428
rect 34495 36097 45047 36393
rect 45423 36097 45430 36393
rect 34495 36060 45430 36097
rect 53690 36368 54350 36390
rect 34495 36052 45110 36060
rect 34240 36020 45110 36052
rect 53690 36025 53712 36368
rect 53625 35672 53712 36025
rect 54328 36025 54350 36368
rect 56340 36130 57080 36600
rect 58440 36160 59180 36600
rect 58725 36145 58940 36160
rect 60540 36070 61280 36600
rect 62640 36090 63380 36600
rect 54328 35672 54895 36025
rect 53625 35585 54895 35672
rect 33900 33138 34000 33145
rect 33900 33125 33924 33138
rect 33455 33086 33924 33125
rect 33976 33125 34000 33138
rect 33976 33093 34520 33125
rect 33976 33086 34244 33093
rect 33455 32988 34244 33086
rect 33455 32936 33601 32988
rect 33653 32936 33856 32988
rect 33908 32957 34244 32988
rect 34460 32957 34520 33093
rect 33908 32936 34520 32957
rect 33455 32925 34520 32936
rect 53710 33050 54520 35585
rect 33045 32863 33910 32875
rect 33045 32811 33466 32863
rect 33518 32811 33726 32863
rect 33778 32811 33910 32863
rect 33045 32743 33910 32811
rect 33045 32691 33796 32743
rect 33848 32691 33910 32743
rect 33045 32675 33910 32691
rect 53710 32715 55650 33050
rect 53710 32240 55996 32715
rect 55432 32200 55996 32240
rect 33260 32128 33380 32155
rect 33260 32076 33294 32128
rect 33346 32076 33380 32128
rect 33260 32064 33380 32076
rect 33260 32012 33294 32064
rect 33346 32012 33380 32064
rect 33260 31990 33380 32012
rect 52150 31529 52240 31560
rect 52150 31477 52169 31529
rect 52221 31477 52240 31529
rect 52150 31465 52240 31477
rect 52150 31413 52169 31465
rect 52221 31413 52240 31465
rect 52150 31401 52240 31413
rect 52150 31349 52169 31401
rect 52221 31349 52240 31401
rect 52150 31337 52240 31349
rect 52150 31285 52169 31337
rect 52221 31285 52240 31337
rect 52150 31273 52240 31285
rect 52150 31221 52169 31273
rect 52221 31221 52240 31273
rect 36440 31178 36900 31200
rect 52150 31190 52240 31221
rect 54804 31529 55168 31558
rect 54804 31233 54838 31529
rect 55134 31233 55168 31529
rect 54804 31204 55168 31233
rect 36440 31122 36482 31178
rect 36538 31176 36562 31178
rect 36618 31176 36642 31178
rect 36698 31176 36722 31178
rect 36778 31176 36802 31178
rect 36538 31124 36548 31176
rect 36792 31124 36802 31176
rect 36538 31122 36562 31124
rect 36618 31122 36642 31124
rect 36698 31122 36722 31124
rect 36778 31122 36802 31124
rect 36858 31122 36900 31178
rect 36440 31100 36900 31122
rect 35740 30959 35980 31000
rect 35740 30651 35770 30959
rect 35950 30651 35980 30959
rect 35740 30610 35980 30651
rect 35760 27001 45180 27030
rect 35760 26949 35785 27001
rect 35837 26949 45180 27001
rect 35760 26937 45180 26949
rect 35760 26885 35785 26937
rect 35837 26885 45180 26937
rect 35760 26873 45180 26885
rect 35760 26821 35785 26873
rect 35837 26821 45180 26873
rect 35760 26809 45180 26821
rect 35760 26757 35785 26809
rect 35837 26757 45180 26809
rect 35760 26745 45180 26757
rect 35760 26693 35785 26745
rect 35837 26693 45180 26745
rect 35760 26681 45180 26693
rect 35760 26629 35785 26681
rect 35837 26629 45180 26681
rect 35760 26600 45180 26629
rect 52145 26438 52235 26440
rect 52145 26386 52164 26438
rect 52216 26386 52235 26438
rect 54882 26420 55210 26422
rect 52145 26374 52235 26386
rect 52145 26322 52164 26374
rect 52216 26322 52235 26374
rect 52145 26310 52235 26322
rect 52145 26258 52164 26310
rect 52216 26258 52235 26310
rect 52145 26246 52235 26258
rect 52145 26194 52164 26246
rect 52216 26194 52235 26246
rect 52145 26182 52235 26194
rect 52145 26130 52164 26182
rect 52216 26130 52235 26182
rect 52145 26118 52235 26130
rect 52145 26066 52164 26118
rect 52216 26066 52235 26118
rect 54840 26404 55210 26420
rect 54840 26108 54877 26404
rect 55173 26108 55210 26404
rect 54840 26090 55210 26108
rect 52145 26065 52235 26066
rect 36420 25538 36940 25560
rect 36420 25536 36452 25538
rect 36508 25536 36532 25538
rect 36588 25536 36612 25538
rect 36668 25536 36692 25538
rect 36748 25536 36772 25538
rect 36828 25536 36852 25538
rect 36908 25536 36940 25538
rect 36420 25484 36430 25536
rect 36610 25484 36612 25536
rect 36674 25484 36686 25536
rect 36748 25484 36750 25536
rect 36930 25484 36940 25536
rect 36420 25482 36452 25484
rect 36508 25482 36532 25484
rect 36588 25482 36612 25484
rect 36668 25482 36692 25484
rect 36748 25482 36772 25484
rect 36828 25482 36852 25484
rect 36908 25482 36940 25484
rect 36420 25470 36940 25482
rect 34665 25304 36160 25345
rect 34665 25252 36074 25304
rect 36126 25252 36160 25304
rect 34665 25240 36160 25252
rect 34665 25188 36074 25240
rect 36126 25188 36160 25240
rect 34665 25176 36160 25188
rect 34665 25124 36074 25176
rect 36126 25124 36160 25176
rect 34665 25112 36160 25124
rect 34665 25060 36074 25112
rect 36126 25060 36160 25112
rect 34665 25020 36160 25060
rect 53900 24570 55890 25380
rect 32940 24448 33300 24465
rect 32940 24396 32966 24448
rect 33018 24396 33030 24448
rect 33082 24396 33094 24448
rect 33146 24396 33158 24448
rect 33210 24396 33222 24448
rect 33274 24396 33300 24448
rect 32940 24380 33300 24396
rect 53900 22045 54710 24570
rect 53600 21958 54895 22045
rect 53600 21605 53717 21958
rect 53680 21262 53717 21605
rect 54573 21605 54895 21958
rect 54573 21262 54610 21605
rect 53680 21230 54610 21262
rect 56340 21035 57080 21530
rect 58440 21035 59180 21550
rect 60540 21035 61280 21540
rect 62895 21440 63110 21475
rect 62640 21035 63380 21440
rect 54785 21030 63380 21035
rect 54780 20993 63380 21030
rect 54780 20537 54832 20993
rect 55208 20840 63380 20993
rect 55208 20537 63370 20840
rect 54780 20430 63370 20537
<< via2 >>
rect 43737 37952 44193 38248
rect 47717 36643 47719 36673
rect 47719 36643 47771 36673
rect 47771 36643 47773 36673
rect 47717 36631 47773 36643
rect 47717 36617 47719 36631
rect 47719 36617 47771 36631
rect 47771 36617 47773 36631
rect 47717 36579 47719 36593
rect 47719 36579 47771 36593
rect 47771 36579 47773 36593
rect 47717 36567 47773 36579
rect 47717 36537 47719 36567
rect 47719 36537 47771 36567
rect 47771 36537 47773 36567
rect 48187 36643 48189 36673
rect 48189 36643 48241 36673
rect 48241 36643 48243 36673
rect 48187 36631 48243 36643
rect 48187 36617 48189 36631
rect 48189 36617 48241 36631
rect 48241 36617 48243 36631
rect 54812 36622 55188 37158
rect 48187 36579 48189 36593
rect 48189 36579 48241 36593
rect 48241 36579 48243 36593
rect 48187 36567 48243 36579
rect 48187 36537 48189 36567
rect 48189 36537 48241 36567
rect 48241 36537 48243 36567
rect 34279 36052 34495 36428
rect 45047 36097 45423 36393
rect 53712 35672 54328 36368
rect 34244 32957 34460 33093
rect 54838 31233 55134 31529
rect 36482 31176 36538 31178
rect 36562 31176 36618 31178
rect 36642 31176 36698 31178
rect 36722 31176 36778 31178
rect 36802 31176 36858 31178
rect 36482 31124 36484 31176
rect 36484 31124 36536 31176
rect 36536 31124 36538 31176
rect 36562 31124 36600 31176
rect 36600 31124 36612 31176
rect 36612 31124 36618 31176
rect 36642 31124 36664 31176
rect 36664 31124 36676 31176
rect 36676 31124 36698 31176
rect 36722 31124 36728 31176
rect 36728 31124 36740 31176
rect 36740 31124 36778 31176
rect 36802 31124 36804 31176
rect 36804 31124 36856 31176
rect 36856 31124 36858 31176
rect 36482 31122 36538 31124
rect 36562 31122 36618 31124
rect 36642 31122 36698 31124
rect 36722 31122 36778 31124
rect 36802 31122 36858 31124
rect 35792 30657 35928 30953
rect 54877 26108 55173 26404
rect 36452 25536 36508 25538
rect 36532 25536 36588 25538
rect 36612 25536 36668 25538
rect 36692 25536 36748 25538
rect 36772 25536 36828 25538
rect 36852 25536 36908 25538
rect 36452 25484 36482 25536
rect 36482 25484 36494 25536
rect 36494 25484 36508 25536
rect 36532 25484 36546 25536
rect 36546 25484 36558 25536
rect 36558 25484 36588 25536
rect 36612 25484 36622 25536
rect 36622 25484 36668 25536
rect 36692 25484 36738 25536
rect 36738 25484 36748 25536
rect 36772 25484 36802 25536
rect 36802 25484 36814 25536
rect 36814 25484 36828 25536
rect 36852 25484 36866 25536
rect 36866 25484 36878 25536
rect 36878 25484 36908 25536
rect 36452 25482 36508 25484
rect 36532 25482 36588 25484
rect 36612 25482 36668 25484
rect 36692 25482 36748 25484
rect 36772 25482 36828 25484
rect 36852 25482 36908 25484
rect 53717 21262 54573 21958
rect 54832 20537 55208 20993
<< metal3 >>
rect 43670 38248 44270 38310
rect 43670 37952 43737 38248
rect 44193 37952 44270 38248
rect 34190 36428 34635 36460
rect 34190 36397 34279 36428
rect 34495 36397 34635 36428
rect 34190 36093 34258 36397
rect 34562 36093 34635 36397
rect 34190 36052 34279 36093
rect 34495 36052 34635 36093
rect 34190 36020 34635 36052
rect 34190 33093 34540 36020
rect 34190 32957 34244 33093
rect 34460 32957 34540 33093
rect 34190 32330 34540 32957
rect 34240 32200 34540 32330
rect 36410 32470 36940 32500
rect 43670 32470 44270 37952
rect 45000 36397 45470 38130
rect 54790 37158 55250 37200
rect 54790 36795 54812 37158
rect 47220 36673 47790 36710
rect 47220 36617 47717 36673
rect 47773 36617 47790 36673
rect 47220 36593 47790 36617
rect 47220 36537 47717 36593
rect 47773 36537 47790 36593
rect 47220 36500 47790 36537
rect 48170 36673 49720 36710
rect 48170 36617 48187 36673
rect 48243 36617 49720 36673
rect 48170 36593 49720 36617
rect 48170 36537 48187 36593
rect 48243 36537 49720 36593
rect 48170 36500 49720 36537
rect 54785 36622 54812 36795
rect 55188 36622 55250 37158
rect 45000 36093 45043 36397
rect 45427 36093 45470 36397
rect 45000 36020 45470 36093
rect 53612 36372 54420 36468
rect 53612 35668 53708 36372
rect 54332 35668 54420 36372
rect 53612 35578 54420 35668
rect 54785 36083 54858 36622
rect 55162 36083 55250 36622
rect 56840 37142 57650 37800
rect 56840 36678 56978 37142
rect 57522 36678 57650 37142
rect 56840 36590 57650 36678
rect 36410 32422 44270 32470
rect 36410 31958 36488 32422
rect 36872 31958 44270 32422
rect 36410 31880 44270 31958
rect 36410 31320 36940 31880
rect 54785 31578 55250 36083
rect 54785 31576 56340 31578
rect 54782 31529 56340 31576
rect 54782 31233 54838 31529
rect 55134 31233 56340 31529
rect 36440 31178 36900 31200
rect 36440 31122 36482 31178
rect 36538 31122 36562 31178
rect 36618 31122 36642 31178
rect 36698 31122 36722 31178
rect 36778 31122 36802 31178
rect 36858 31122 36900 31178
rect 54782 31176 56340 31233
rect 36440 31100 36900 31122
rect 35740 30957 35980 31000
rect 35740 30653 35788 30957
rect 35932 30653 35980 30957
rect 35740 30610 35980 30653
rect 57735 30242 58240 30245
rect 55465 30199 55925 30220
rect 55465 29895 55503 30199
rect 55887 29895 55925 30199
rect 55465 29875 55925 29895
rect 57480 29855 57720 30020
rect 57735 29858 57755 30242
rect 58219 29858 58240 30242
rect 61085 30194 62590 30270
rect 57735 29855 58240 29858
rect 59610 30057 59755 30060
rect 59300 29673 59610 29800
rect 59754 29800 59755 30057
rect 61085 29810 61875 30194
rect 62499 29810 62590 30194
rect 59754 29673 59780 29800
rect 61085 29785 62590 29810
rect 59300 29490 59780 29673
rect 59620 28109 59860 28120
rect 56407 27820 56420 28090
rect 55650 27750 55670 27770
rect 57710 27764 58235 27765
rect 55465 27719 55950 27750
rect 55465 27415 55475 27719
rect 55939 27415 55950 27719
rect 55465 27385 55950 27415
rect 57710 27380 57740 27764
rect 58204 27380 58235 27764
rect 59620 27565 59628 28109
rect 59852 27565 59860 28109
rect 59620 27555 59860 27565
rect 61090 27784 62625 27835
rect 61090 27400 61868 27784
rect 62572 27400 62625 27784
rect 61090 27360 62625 27400
rect 54790 26456 55260 26460
rect 54790 26407 56470 26456
rect 54790 26103 54868 26407
rect 55172 26404 56470 26407
rect 55173 26108 56470 26404
rect 55172 26103 56470 26108
rect 54790 26060 56470 26103
rect 54795 26054 56470 26060
rect 36430 25538 36930 25540
rect 36430 25482 36452 25538
rect 36508 25482 36532 25538
rect 36588 25482 36612 25538
rect 36668 25482 36692 25538
rect 36748 25482 36772 25538
rect 36828 25482 36852 25538
rect 36908 25482 36930 25538
rect 36430 25480 36930 25482
rect 33845 24612 36555 24695
rect 33845 24148 34563 24612
rect 35747 24148 36555 24612
rect 33845 24090 36555 24148
rect 54795 23542 55260 26054
rect 54795 22598 54888 23542
rect 55112 22598 55260 23542
rect 53610 21962 54670 22040
rect 53610 21258 53713 21962
rect 54577 21258 54670 21962
rect 53610 21170 54670 21258
rect 54795 20993 55260 22598
rect 54795 20845 54832 20993
rect 54800 20537 54832 20845
rect 55208 20537 55260 20993
rect 54800 20430 55260 20537
<< via3 >>
rect 34258 36093 34279 36397
rect 34279 36093 34495 36397
rect 34495 36093 34562 36397
rect 54858 36622 55162 37107
rect 45043 36393 45427 36397
rect 45043 36097 45047 36393
rect 45047 36097 45423 36393
rect 45423 36097 45427 36393
rect 45043 36093 45427 36097
rect 53708 36368 54332 36372
rect 53708 35672 53712 36368
rect 53712 35672 54328 36368
rect 54328 35672 54332 36368
rect 53708 35668 54332 35672
rect 54858 36083 55162 36622
rect 56978 36678 57522 37142
rect 36488 31958 36872 32422
rect 35788 30953 35932 30957
rect 35788 30657 35792 30953
rect 35792 30657 35928 30953
rect 35928 30657 35932 30953
rect 35788 30653 35932 30657
rect 55503 29895 55887 30199
rect 57755 29858 58219 30242
rect 59610 29673 59754 30057
rect 61875 29810 62499 30194
rect 55475 27415 55939 27719
rect 57740 27380 58204 27764
rect 59628 27565 59852 28109
rect 61868 27400 62572 27784
rect 54868 26404 55172 26407
rect 54868 26108 54877 26404
rect 54877 26108 55172 26404
rect 54868 26103 55172 26108
rect 34563 24148 35747 24612
rect 54888 22598 55112 23542
rect 53713 21958 54577 21962
rect 53713 21262 53717 21958
rect 53717 21262 54573 21958
rect 54573 21262 54577 21958
rect 53713 21258 54577 21262
<< metal4 >>
rect 52260 36470 52850 37560
rect 54780 37142 65400 37240
rect 54780 37107 56978 37142
rect 52260 36468 54190 36470
rect 34190 36397 34630 36460
rect 34190 36093 34258 36397
rect 34562 36093 34630 36397
rect 34190 36020 34630 36093
rect 45000 36397 45470 36460
rect 45000 36093 45043 36397
rect 45427 36093 45470 36397
rect 45000 36030 45470 36093
rect 52260 36372 54420 36468
rect 52260 35860 53708 36372
rect 53612 35668 53708 35860
rect 54332 35668 54420 36372
rect 54780 36083 54858 37107
rect 55162 37028 56978 37107
rect 57522 37028 65400 37142
rect 55162 36792 56972 37028
rect 57528 36792 65400 37028
rect 55162 36678 56978 36792
rect 57522 36678 65400 36792
rect 55162 36600 65400 36678
rect 55162 36083 55250 36600
rect 56840 36590 57650 36600
rect 54780 36000 55250 36083
rect 53612 35578 54420 35668
rect 36410 32422 36940 32500
rect 36410 31958 36488 32422
rect 36872 31958 36940 32422
rect 36410 31840 36940 31958
rect 35740 30957 36320 31000
rect 35740 30653 35788 30957
rect 35932 30653 36320 30957
rect 35740 30610 36320 30653
rect 61810 30300 62585 30475
rect 55435 30199 56170 30260
rect 55435 29895 55503 30199
rect 55887 30193 56170 30199
rect 56040 29957 56170 30193
rect 55887 29895 56170 29957
rect 55435 29850 56170 29895
rect 57695 30242 58260 30270
rect 57695 29858 57755 30242
rect 58219 29858 58260 30242
rect 61810 30194 62167 30300
rect 62403 30194 62585 30300
rect 59865 30158 60165 30190
rect 59865 30095 59902 30158
rect 57695 29835 58260 29858
rect 59600 30057 59902 30095
rect 59600 29673 59610 30057
rect 59754 29922 59902 30057
rect 60138 29922 60165 30158
rect 59754 29895 60165 29922
rect 59754 29673 59775 29895
rect 61810 29810 61875 30194
rect 62499 29810 62585 30194
rect 61810 29780 62585 29810
rect 59600 29655 59775 29673
rect 59600 28109 59885 28140
rect 55440 27719 56175 27820
rect 55440 27415 55475 27719
rect 55939 27665 56175 27719
rect 56035 27429 56175 27665
rect 55939 27415 56175 27429
rect 55440 27355 56175 27415
rect 57695 27764 58255 27790
rect 57695 27380 57740 27764
rect 58204 27380 58255 27764
rect 59600 27565 59628 28109
rect 59852 27735 59885 28109
rect 61810 27784 62620 27830
rect 59852 27713 60200 27735
rect 59852 27565 59924 27713
rect 59600 27510 59924 27565
rect 59885 27477 59924 27510
rect 60160 27477 60200 27713
rect 59885 27465 60200 27477
rect 57695 27360 58255 27380
rect 61810 27400 61868 27784
rect 62572 27598 62620 27784
rect 61810 27362 62019 27400
rect 62255 27362 62339 27400
rect 62575 27362 62620 27598
rect 61810 27225 62620 27362
rect 54790 26407 55250 26460
rect 54790 26103 54868 26407
rect 55172 26103 55250 26407
rect 54790 26060 55250 26103
rect 34440 24612 35960 24700
rect 34440 24498 34563 24612
rect 35747 24498 35960 24612
rect 34440 24262 34557 24498
rect 35753 24262 35960 24498
rect 34440 24148 34563 24262
rect 35747 24148 35960 24262
rect 34440 23320 35960 24148
rect 54760 23542 55240 23630
rect 54760 23508 54888 23542
rect 55112 23508 55240 23542
rect 54760 23272 54882 23508
rect 55118 23272 55240 23508
rect 54760 23188 54888 23272
rect 55112 23188 55240 23272
rect 54760 22952 54882 23188
rect 55118 22952 55240 23188
rect 54760 22868 54888 22952
rect 55112 22868 55240 22952
rect 54760 22632 54882 22868
rect 55118 22632 55240 22868
rect 54760 22598 54888 22632
rect 55112 22598 55240 22632
rect 54760 22520 55240 22598
rect 53610 21962 54670 22040
rect 53610 21888 53713 21962
rect 54577 21888 54670 21962
rect 53610 21332 53707 21888
rect 54583 21332 54670 21888
rect 53610 21258 53713 21332
rect 54577 21258 54670 21332
rect 53610 21170 54670 21258
<< via4 >>
rect 34292 36127 34528 36363
rect 45117 36127 45353 36363
rect 53742 35742 54298 36298
rect 54892 36797 55128 37033
rect 56972 36792 56978 37028
rect 56978 36792 57208 37028
rect 57292 36792 57522 37028
rect 57522 36792 57528 37028
rect 54892 36477 55128 36713
rect 54892 36157 55128 36393
rect 36562 32072 36798 32308
rect 55804 29957 55887 30193
rect 55887 29957 56040 30193
rect 57869 29937 58105 30173
rect 62167 30194 62403 30300
rect 59902 29922 60138 30158
rect 62167 30064 62403 30194
rect 55799 27429 55939 27665
rect 55939 27429 56035 27665
rect 57857 27457 58093 27693
rect 59924 27477 60160 27713
rect 62019 27400 62255 27598
rect 62339 27400 62572 27598
rect 62572 27400 62575 27598
rect 62019 27362 62255 27400
rect 62339 27362 62575 27400
rect 54902 26137 55138 26373
rect 34557 24262 34563 24498
rect 34563 24262 34793 24498
rect 34877 24262 35113 24498
rect 35197 24262 35433 24498
rect 35517 24262 35747 24498
rect 35747 24262 35753 24498
rect 54882 23272 54888 23508
rect 54888 23272 55112 23508
rect 55112 23272 55118 23508
rect 54882 22952 54888 23188
rect 54888 22952 55112 23188
rect 55112 22952 55118 23188
rect 54882 22632 54888 22868
rect 54888 22632 55112 22868
rect 55112 22632 55118 22868
rect 53707 21332 53713 21888
rect 53713 21332 54577 21888
rect 54577 21332 54583 21888
<< metal5 >>
rect 54780 37033 57650 37240
rect 54780 36797 54892 37033
rect 55128 37028 57650 37033
rect 55128 36797 56972 37028
rect 54780 36792 56972 36797
rect 57208 36792 57292 37028
rect 57528 36792 57650 37028
rect 54780 36713 57650 36792
rect 54780 36477 54892 36713
rect 55128 36590 57650 36713
rect 55128 36477 55330 36590
rect 53612 36460 54420 36468
rect 34170 36363 54420 36460
rect 34170 36127 34292 36363
rect 34528 36127 45117 36363
rect 45353 36298 54420 36363
rect 45353 36127 53742 36298
rect 34170 35742 53742 36127
rect 54298 35742 54420 36298
rect 34170 35640 54420 35742
rect 53612 35578 54420 35640
rect 54780 36393 55330 36477
rect 54780 36157 54892 36393
rect 55128 36157 55330 36393
rect 36330 32308 37030 32510
rect 36330 32072 36562 32308
rect 36798 32072 37030 32308
rect 36330 24710 37030 32072
rect 34480 24498 37040 24710
rect 34480 24262 34557 24498
rect 34793 24262 34877 24498
rect 35113 24262 35197 24498
rect 35433 24262 35517 24498
rect 35753 24262 37040 24498
rect 34480 24080 37040 24262
rect 53630 22040 54080 35578
rect 54780 35180 55330 36157
rect 54550 34620 55330 35180
rect 54550 26373 55250 34620
rect 62015 30300 62555 30435
rect 55705 30193 56135 30230
rect 55705 29957 55804 30193
rect 56040 29957 56135 30193
rect 55705 29920 56135 29957
rect 57695 30173 58260 30270
rect 57695 29937 57869 30173
rect 58105 29937 58260 30173
rect 57695 29910 58260 29937
rect 59865 30190 59895 30215
rect 59865 30158 60165 30190
rect 59865 29922 59902 30158
rect 60138 29922 60165 30158
rect 62015 30064 62167 30300
rect 62403 30064 62555 30300
rect 62015 29930 62555 30064
rect 57695 29835 58265 29910
rect 59865 29895 60165 29922
rect 55710 27665 56125 27705
rect 55710 27429 55799 27665
rect 56035 27429 56125 27665
rect 55710 27390 56125 27429
rect 57685 27693 58260 27790
rect 57685 27457 57857 27693
rect 58093 27457 58260 27693
rect 57685 27360 58260 27457
rect 59875 27713 60200 27740
rect 59875 27477 59924 27713
rect 60160 27477 60200 27713
rect 59875 27400 60200 27477
rect 62015 27598 62580 27700
rect 62015 27362 62019 27598
rect 62255 27362 62339 27598
rect 62575 27362 62580 27598
rect 62015 27260 62580 27362
rect 54550 26137 54902 26373
rect 55138 26137 55250 26373
rect 54550 23508 55250 26137
rect 54550 23272 54882 23508
rect 55118 23272 55250 23508
rect 54550 23188 55250 23272
rect 54550 22952 54882 23188
rect 55118 22952 55250 23188
rect 54550 22868 55250 22952
rect 54550 22632 54882 22868
rect 55118 22632 55250 22868
rect 54550 22520 55250 22632
rect 53610 21888 54670 22040
rect 53610 21332 53707 21888
rect 54583 21332 54670 21888
rect 53610 21170 54670 21332
use core_osc  X1
timestamp 1663011646
transform 1 0 46065 0 1 21045
box 9175 3425 16085 12111
use buffer_amp_vop  X3
timestamp 1663011646
transform 1 0 26070 0 1 10600
box 10225 10400 29180 26030
use cap_bank  X4
timestamp 1663011646
transform 1 0 52305 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X5
timestamp 1663011646
transform 1 0 54405 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X6
timestamp 1663011646
transform 1 0 52305 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X7
timestamp 1663011646
transform 1 0 54405 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X8
timestamp 1663011646
transform 1 0 56505 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X9
timestamp 1663011646
transform 1 0 58605 0 1 22905
box 3300 -1540 5112 5514
use cap_bank  X10
timestamp 1663011646
transform 1 0 56505 0 -1 34725
box 3300 -1540 5112 5514
use cap_bank  X11
timestamp 1663011646
transform 1 0 58605 0 -1 34725
box 3300 -1540 5112 5514
use bias_calc  bias_calc_0
timestamp 1663011646
transform 1 0 14295 0 1 25060
box 16856 -965 21340 7275
use output_buffer  output_buffer_0
timestamp 1663011646
transform 1 0 34825 0 1 39195
box 8845 -1865 22825 2475
use sky130_fd_pr__pfet_01v8_lvt_75KH85  sky130_fd_pr__pfet_01v8_lvt_75KH85_0
timestamp 1663011646
transform 1 0 33689 0 1 32864
box -359 -284 359 284
<< labels >>
rlabel metal5 s 53630 21190 54080 36450 4 VDD
port 1 nsew
rlabel metal5 s 36330 24100 37030 32510 4 GND
port 2 nsew
rlabel metal1 s 64850 21365 64910 36265 4 CTRL1
port 3 nsew
rlabel metal1 s 64595 21725 64655 35905 4 CTRL2
port 4 nsew
rlabel metal1 s 64345 22265 64405 35365 4 CTRL3
port 5 nsew
rlabel metal1 s 64080 22855 64140 34775 4 CTRL4
port 6 nsew
rlabel metal1 s 63845 23765 63905 33865 4 CTRL5
port 7 nsew
rlabel metal2 s 60540 36070 61280 37200 4 GND
port 2 nsew
<< end >>
