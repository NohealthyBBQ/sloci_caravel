magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -173 172 -115 178
rect 19 172 77 178
rect 211 172 269 178
rect -173 138 -161 172
rect 19 138 31 172
rect 211 138 223 172
rect -173 132 -115 138
rect 19 132 77 138
rect 211 132 269 138
rect -269 -138 -211 -132
rect -77 -138 -19 -132
rect 115 -138 173 -132
rect -269 -172 -257 -138
rect -77 -172 -65 -138
rect 115 -172 127 -138
rect -269 -178 -211 -172
rect -77 -178 -19 -172
rect 115 -178 173 -172
<< pwell >>
rect -445 -300 445 300
<< nmoslvt >>
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
<< ndiff >>
rect -317 85 -255 100
rect -317 51 -305 85
rect -271 51 -255 85
rect -317 17 -255 51
rect -317 -17 -305 17
rect -271 -17 -255 17
rect -317 -51 -255 -17
rect -317 -85 -305 -51
rect -271 -85 -255 -51
rect -317 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 317 100
rect 255 51 271 85
rect 305 51 317 85
rect 255 17 317 51
rect 255 -17 271 17
rect 305 -17 317 17
rect 255 -51 317 -17
rect 255 -85 271 -51
rect 305 -85 317 -51
rect 255 -100 317 -85
<< ndiffc >>
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
<< psubdiff >>
rect -419 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 419 274
rect -419 153 -385 240
rect -419 85 -385 119
rect 385 153 419 240
rect -419 17 -385 51
rect -419 -51 -385 -17
rect -419 -119 -385 -85
rect 385 85 419 119
rect 385 17 419 51
rect 385 -51 419 -17
rect -419 -240 -385 -153
rect 385 -119 419 -85
rect 385 -240 419 -153
rect -419 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 419 -240
<< psubdiffcont >>
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect -419 119 -385 153
rect 385 119 419 153
rect -419 51 -385 85
rect -419 -17 -385 17
rect -419 -85 -385 -51
rect 385 51 419 85
rect 385 -17 419 17
rect 385 -85 419 -51
rect -419 -153 -385 -119
rect 385 -153 419 -119
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
<< poly >>
rect -177 172 -111 188
rect -177 138 -161 172
rect -127 138 -111 172
rect -255 100 -225 126
rect -177 122 -111 138
rect 15 172 81 188
rect 15 138 31 172
rect 65 138 81 172
rect -159 100 -129 122
rect -63 100 -33 126
rect 15 122 81 138
rect 207 172 273 188
rect 207 138 223 172
rect 257 138 273 172
rect 33 100 63 122
rect 129 100 159 126
rect 207 122 273 138
rect 225 100 255 122
rect -255 -122 -225 -100
rect -273 -138 -207 -122
rect -159 -126 -129 -100
rect -63 -122 -33 -100
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -273 -188 -207 -172
rect -81 -138 -15 -122
rect 33 -126 63 -100
rect 129 -122 159 -100
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect -81 -188 -15 -172
rect 111 -138 177 -122
rect 225 -126 255 -100
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 111 -188 177 -172
<< polycont >>
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
<< locali >>
rect -419 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 419 274
rect -419 153 -385 240
rect -177 138 -161 172
rect -127 138 -111 172
rect 15 138 31 172
rect 65 138 81 172
rect 207 138 223 172
rect 257 138 273 172
rect 385 153 419 240
rect -419 85 -385 119
rect -419 17 -385 51
rect -419 -51 -385 -17
rect -419 -119 -385 -85
rect -305 85 -271 104
rect -305 17 -271 19
rect -305 -19 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 19
rect 271 -19 305 -17
rect 271 -104 305 -85
rect 385 85 419 119
rect 385 17 419 51
rect 385 -51 419 -17
rect 385 -119 419 -85
rect -419 -240 -385 -153
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 385 -240 419 -153
rect -419 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 419 -240
<< viali >>
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
<< metal1 >>
rect -173 172 -115 178
rect -173 138 -161 172
rect -127 138 -115 172
rect -173 132 -115 138
rect 19 172 77 178
rect 19 138 31 172
rect 65 138 77 172
rect 19 132 77 138
rect 211 172 269 178
rect 211 138 223 172
rect 257 138 269 172
rect 211 132 269 138
rect -311 53 -265 100
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -100 -265 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 265 53 311 100
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -100 311 -53
rect -269 -138 -211 -132
rect -269 -172 -257 -138
rect -223 -172 -211 -138
rect -269 -178 -211 -172
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -31 -172 -19 -138
rect -77 -178 -19 -172
rect 115 -138 173 -132
rect 115 -172 127 -138
rect 161 -172 173 -138
rect 115 -178 173 -172
<< properties >>
string FIXED_BBOX -402 -257 402 257
<< end >>
