magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -700 -500 2900 3100
<< nsubdiff >>
rect -500 2967 2700 3000
rect -500 2933 827 2967
rect 861 2933 895 2967
rect 929 2933 963 2967
rect 997 2933 1031 2967
rect 1065 2933 1099 2967
rect 1133 2933 1167 2967
rect 1201 2933 1235 2967
rect 1269 2933 1303 2967
rect 1337 2933 1371 2967
rect 1405 2933 1439 2967
rect 1473 2933 2700 2967
rect -500 2900 2700 2933
rect -500 1691 -400 2900
rect -500 1657 -467 1691
rect -433 1657 -400 1691
rect -500 1623 -400 1657
rect -500 1589 -467 1623
rect -433 1589 -400 1623
rect -500 1555 -400 1589
rect -500 1521 -467 1555
rect -433 1521 -400 1555
rect -500 1487 -400 1521
rect -500 1453 -467 1487
rect -433 1453 -400 1487
rect -500 1419 -400 1453
rect -500 1385 -467 1419
rect -433 1385 -400 1419
rect -500 1351 -400 1385
rect -500 1317 -467 1351
rect -433 1317 -400 1351
rect -500 1283 -400 1317
rect -500 1249 -467 1283
rect -433 1249 -400 1283
rect -500 1215 -400 1249
rect -500 1181 -467 1215
rect -433 1181 -400 1215
rect -500 1147 -400 1181
rect -500 1113 -467 1147
rect -433 1113 -400 1147
rect -500 1079 -400 1113
rect -500 1045 -467 1079
rect -433 1045 -400 1079
rect -500 1011 -400 1045
rect -500 977 -467 1011
rect -433 977 -400 1011
rect -500 943 -400 977
rect -500 909 -467 943
rect -433 909 -400 943
rect -500 -300 -400 909
rect 2600 1691 2700 2900
rect 2600 1657 2633 1691
rect 2667 1657 2700 1691
rect 2600 1623 2700 1657
rect 2600 1589 2633 1623
rect 2667 1589 2700 1623
rect 2600 1555 2700 1589
rect 2600 1521 2633 1555
rect 2667 1521 2700 1555
rect 2600 1487 2700 1521
rect 2600 1453 2633 1487
rect 2667 1453 2700 1487
rect 2600 1419 2700 1453
rect 2600 1385 2633 1419
rect 2667 1385 2700 1419
rect 2600 1351 2700 1385
rect 2600 1317 2633 1351
rect 2667 1317 2700 1351
rect 2600 1283 2700 1317
rect 2600 1249 2633 1283
rect 2667 1249 2700 1283
rect 2600 1215 2700 1249
rect 2600 1181 2633 1215
rect 2667 1181 2700 1215
rect 2600 1147 2700 1181
rect 2600 1113 2633 1147
rect 2667 1113 2700 1147
rect 2600 1079 2700 1113
rect 2600 1045 2633 1079
rect 2667 1045 2700 1079
rect 2600 1011 2700 1045
rect 2600 977 2633 1011
rect 2667 977 2700 1011
rect 2600 943 2700 977
rect 2600 909 2633 943
rect 2667 909 2700 943
rect 2600 -300 2700 909
rect -500 -333 2700 -300
rect -500 -367 827 -333
rect 861 -367 895 -333
rect 929 -367 963 -333
rect 997 -367 1031 -333
rect 1065 -367 1099 -333
rect 1133 -367 1167 -333
rect 1201 -367 1235 -333
rect 1269 -367 1303 -333
rect 1337 -367 1371 -333
rect 1405 -367 1439 -333
rect 1473 -367 2700 -333
rect -500 -400 2700 -367
<< nsubdiffcont >>
rect 827 2933 861 2967
rect 895 2933 929 2967
rect 963 2933 997 2967
rect 1031 2933 1065 2967
rect 1099 2933 1133 2967
rect 1167 2933 1201 2967
rect 1235 2933 1269 2967
rect 1303 2933 1337 2967
rect 1371 2933 1405 2967
rect 1439 2933 1473 2967
rect -467 1657 -433 1691
rect -467 1589 -433 1623
rect -467 1521 -433 1555
rect -467 1453 -433 1487
rect -467 1385 -433 1419
rect -467 1317 -433 1351
rect -467 1249 -433 1283
rect -467 1181 -433 1215
rect -467 1113 -433 1147
rect -467 1045 -433 1079
rect -467 977 -433 1011
rect -467 909 -433 943
rect 2633 1657 2667 1691
rect 2633 1589 2667 1623
rect 2633 1521 2667 1555
rect 2633 1453 2667 1487
rect 2633 1385 2667 1419
rect 2633 1317 2667 1351
rect 2633 1249 2667 1283
rect 2633 1181 2667 1215
rect 2633 1113 2667 1147
rect 2633 1045 2667 1079
rect 2633 977 2667 1011
rect 2633 909 2667 943
rect 827 -367 861 -333
rect 895 -367 929 -333
rect 963 -367 997 -333
rect 1031 -367 1065 -333
rect 1099 -367 1133 -333
rect 1167 -367 1201 -333
rect 1235 -367 1269 -333
rect 1303 -367 1337 -333
rect 1371 -367 1405 -333
rect 1439 -367 1473 -333
<< locali >>
rect -500 2967 2700 3000
rect -500 2933 827 2967
rect 861 2933 895 2967
rect 929 2933 963 2967
rect 997 2933 1031 2967
rect 1065 2933 1099 2967
rect 1133 2933 1167 2967
rect 1201 2933 1235 2967
rect 1269 2933 1303 2967
rect 1337 2933 1371 2967
rect 1405 2933 1439 2967
rect 1473 2933 2700 2967
rect -500 2900 2700 2933
rect -500 1691 -400 2900
rect -500 1657 -467 1691
rect -433 1657 -400 1691
rect -500 1623 -400 1657
rect -500 1589 -467 1623
rect -433 1589 -400 1623
rect -500 1555 -400 1589
rect -500 1521 -467 1555
rect -433 1521 -400 1555
rect -500 1487 -400 1521
rect -500 1453 -467 1487
rect -433 1453 -400 1487
rect -500 1419 -400 1453
rect -500 1385 -467 1419
rect -433 1385 -400 1419
rect -500 1351 -400 1385
rect -500 1317 -467 1351
rect -433 1317 -400 1351
rect -500 1283 -400 1317
rect -500 1249 -467 1283
rect -433 1249 -400 1283
rect -500 1215 -400 1249
rect -500 1181 -467 1215
rect -433 1181 -400 1215
rect -500 1147 -400 1181
rect -500 1113 -467 1147
rect -433 1113 -400 1147
rect -500 1079 -400 1113
rect -500 1045 -467 1079
rect -433 1045 -400 1079
rect -500 1011 -400 1045
rect -500 977 -467 1011
rect -433 977 -400 1011
rect -500 943 -400 977
rect -500 909 -467 943
rect -433 909 -400 943
rect -500 -300 -400 909
rect 2600 1691 2700 2900
rect 2600 1657 2633 1691
rect 2667 1657 2700 1691
rect 2600 1623 2700 1657
rect 2600 1589 2633 1623
rect 2667 1589 2700 1623
rect 2600 1555 2700 1589
rect 2600 1521 2633 1555
rect 2667 1521 2700 1555
rect 2600 1487 2700 1521
rect 2600 1453 2633 1487
rect 2667 1453 2700 1487
rect 2600 1419 2700 1453
rect 2600 1385 2633 1419
rect 2667 1385 2700 1419
rect 2600 1351 2700 1385
rect 2600 1317 2633 1351
rect 2667 1317 2700 1351
rect 2600 1283 2700 1317
rect 2600 1249 2633 1283
rect 2667 1249 2700 1283
rect 2600 1215 2700 1249
rect 2600 1181 2633 1215
rect 2667 1181 2700 1215
rect 2600 1147 2700 1181
rect 2600 1113 2633 1147
rect 2667 1113 2700 1147
rect 2600 1079 2700 1113
rect 2600 1045 2633 1079
rect 2667 1045 2700 1079
rect 2600 1011 2700 1045
rect 2600 977 2633 1011
rect 2667 977 2700 1011
rect 2600 943 2700 977
rect 2600 909 2633 943
rect 2667 909 2700 943
rect 2600 -300 2700 909
rect -500 -333 2700 -300
rect -500 -367 827 -333
rect 861 -367 895 -333
rect 929 -367 963 -333
rect 997 -367 1031 -333
rect 1065 -367 1099 -333
rect 1133 -367 1167 -333
rect 1201 -367 1235 -333
rect 1269 -367 1303 -333
rect 1337 -367 1371 -333
rect 1405 -367 1439 -333
rect 1473 -367 2700 -333
rect -500 -400 2700 -367
<< metal1 >>
rect 790 2496 870 2500
rect 790 2444 804 2496
rect 856 2444 870 2496
rect 790 2440 870 2444
rect 1830 2496 1910 2500
rect 1830 2444 1844 2496
rect 1896 2444 1910 2496
rect 1830 2440 1910 2444
rect 30 2416 110 2420
rect 30 2364 44 2416
rect 96 2364 110 2416
rect 30 2360 110 2364
rect 550 2416 630 2420
rect 550 2364 564 2416
rect 616 2364 630 2416
rect 550 2360 630 2364
rect 1050 2416 1130 2420
rect 1050 2364 1064 2416
rect 1116 2364 1130 2416
rect 1050 2360 1130 2364
rect 1570 2416 1650 2420
rect 1570 2364 1584 2416
rect 1636 2364 1650 2416
rect 1570 2360 1650 2364
rect 2090 2416 2170 2420
rect 2090 2364 2104 2416
rect 2156 2364 2170 2416
rect 2090 2360 2170 2364
rect 290 2356 370 2360
rect 290 2304 304 2356
rect 356 2304 370 2356
rect 290 2300 370 2304
rect 1310 2356 1390 2360
rect 1310 2304 1324 2356
rect 1376 2304 1390 2356
rect 1310 2300 1390 2304
rect 98 2202 2096 2250
rect 790 2116 870 2120
rect 790 2064 804 2116
rect 856 2064 870 2116
rect 790 2060 870 2064
rect 1830 2116 1910 2120
rect 1830 2064 1844 2116
rect 1896 2064 1910 2116
rect 1830 2060 1910 2064
rect 30 2056 110 2060
rect 30 2004 44 2056
rect 96 2004 110 2056
rect 30 2000 110 2004
rect 550 2056 630 2060
rect 550 2004 564 2056
rect 616 2004 630 2056
rect 550 2000 630 2004
rect 1050 2056 1130 2060
rect 1050 2004 1064 2056
rect 1116 2004 1130 2056
rect 1050 2000 1130 2004
rect 1570 2056 1650 2060
rect 1570 2004 1584 2056
rect 1636 2004 1650 2056
rect 1570 2000 1650 2004
rect 290 1976 370 1980
rect 290 1924 304 1976
rect 356 1924 370 1976
rect 290 1920 370 1924
rect 1310 1976 1390 1980
rect 1310 1924 1324 1976
rect 1376 1924 1390 1976
rect 1310 1920 1390 1924
rect 1980 1884 2020 2202
rect 2090 2056 2170 2060
rect 2090 2004 2104 2056
rect 2156 2004 2170 2056
rect 2090 2000 2170 2004
rect 98 1838 2096 1884
rect 790 1756 870 1760
rect 790 1704 804 1756
rect 856 1704 870 1756
rect 790 1700 870 1704
rect 1830 1756 1910 1760
rect 1830 1704 1844 1756
rect 1896 1704 1910 1756
rect 1830 1700 1910 1704
rect 30 1696 110 1700
rect 30 1644 44 1696
rect 96 1644 110 1696
rect 30 1640 110 1644
rect 550 1696 630 1700
rect 550 1644 564 1696
rect 616 1644 630 1696
rect 550 1640 630 1644
rect 1050 1696 1130 1700
rect 1050 1644 1064 1696
rect 1116 1644 1130 1696
rect 1050 1640 1130 1644
rect 1570 1696 1650 1700
rect 1570 1644 1584 1696
rect 1636 1644 1650 1696
rect 1570 1640 1650 1644
rect 290 1616 370 1620
rect 290 1564 304 1616
rect 356 1564 370 1616
rect 290 1560 370 1564
rect 1310 1616 1390 1620
rect 1310 1564 1324 1616
rect 1376 1564 1390 1616
rect 1310 1560 1390 1564
rect 1980 1520 2020 1838
rect 2090 1696 2170 1700
rect 2090 1644 2104 1696
rect 2156 1644 2170 1696
rect 2090 1640 2170 1644
rect 98 1472 2096 1520
rect 810 1396 890 1400
rect 810 1344 824 1396
rect 876 1344 890 1396
rect 810 1340 890 1344
rect 1830 1396 1910 1400
rect 1830 1344 1844 1396
rect 1896 1344 1910 1396
rect 1830 1340 1910 1344
rect 30 1336 110 1340
rect 30 1284 44 1336
rect 96 1284 110 1336
rect 30 1280 110 1284
rect 550 1336 630 1340
rect 550 1284 564 1336
rect 616 1284 630 1336
rect 550 1280 630 1284
rect 1050 1336 1130 1340
rect 1050 1284 1064 1336
rect 1116 1284 1130 1336
rect 1050 1280 1130 1284
rect 1570 1336 1650 1340
rect 1570 1284 1584 1336
rect 1636 1284 1650 1336
rect 1570 1280 1650 1284
rect 290 1256 370 1260
rect 290 1204 304 1256
rect 356 1204 370 1256
rect 290 1200 370 1204
rect 1330 1256 1410 1260
rect 1330 1204 1344 1256
rect 1396 1204 1410 1256
rect 1330 1200 1410 1204
rect 1980 1154 2020 1472
rect 2090 1336 2170 1340
rect 2090 1284 2104 1336
rect 2156 1284 2170 1336
rect 2090 1280 2170 1284
rect 98 1108 2096 1154
rect 790 1036 870 1040
rect 790 984 804 1036
rect 856 984 870 1036
rect 790 980 870 984
rect 1830 1036 1910 1040
rect 1830 984 1844 1036
rect 1896 984 1910 1036
rect 1830 980 1910 984
rect 30 956 110 960
rect 30 904 44 956
rect 96 904 110 956
rect 30 900 110 904
rect 550 956 630 960
rect 550 904 564 956
rect 616 904 630 956
rect 550 900 630 904
rect 1050 956 1130 960
rect 1050 904 1064 956
rect 1116 904 1130 956
rect 1050 900 1130 904
rect 1570 956 1650 960
rect 1570 904 1584 956
rect 1636 904 1650 956
rect 1570 900 1650 904
rect 290 896 370 900
rect 290 844 304 896
rect 356 844 370 896
rect 290 840 370 844
rect 1310 896 1390 900
rect 1310 844 1324 896
rect 1376 844 1390 896
rect 1310 840 1390 844
rect 1980 790 2020 1108
rect 2090 956 2170 960
rect 2090 904 2104 956
rect 2156 904 2170 956
rect 2090 900 2170 904
rect 98 742 2096 790
rect 790 656 870 660
rect 790 604 804 656
rect 856 604 870 656
rect 790 600 870 604
rect 1830 656 1910 660
rect 1830 604 1844 656
rect 1896 604 1910 656
rect 1830 600 1910 604
rect 30 596 110 600
rect 30 544 44 596
rect 96 544 110 596
rect 30 540 110 544
rect 550 596 630 600
rect 550 544 564 596
rect 616 544 630 596
rect 550 540 630 544
rect 1050 596 1130 600
rect 1050 544 1064 596
rect 1116 544 1130 596
rect 1050 540 1130 544
rect 1570 596 1650 600
rect 1570 544 1584 596
rect 1636 544 1650 596
rect 1570 540 1650 544
rect 290 516 370 520
rect 290 464 304 516
rect 356 464 370 516
rect 290 460 370 464
rect 1310 516 1390 520
rect 1310 464 1324 516
rect 1376 464 1390 516
rect 1310 460 1390 464
rect 1980 424 2020 742
rect 2090 596 2170 600
rect 2090 544 2104 596
rect 2156 544 2170 596
rect 2090 540 2170 544
rect 98 378 2096 424
rect 790 296 870 300
rect 790 244 804 296
rect 856 244 870 296
rect 790 240 870 244
rect 1830 296 1910 300
rect 1830 244 1844 296
rect 1896 244 1910 296
rect 1830 240 1910 244
rect 30 236 110 240
rect 30 184 44 236
rect 96 184 110 236
rect 30 180 110 184
rect 550 236 630 240
rect 550 184 564 236
rect 616 184 630 236
rect 550 180 630 184
rect 1050 236 1130 240
rect 1050 184 1064 236
rect 1116 184 1130 236
rect 1050 180 1130 184
rect 1570 236 1650 240
rect 1570 184 1584 236
rect 1636 184 1650 236
rect 1570 180 1650 184
rect 290 156 370 160
rect 290 104 304 156
rect 356 104 370 156
rect 290 100 370 104
rect 1310 156 1390 160
rect 1310 104 1324 156
rect 1376 104 1390 156
rect 1310 100 1390 104
rect 1980 60 2020 378
rect 2090 236 2170 240
rect 2090 184 2104 236
rect 2156 184 2170 236
rect 2090 180 2170 184
rect 98 12 2096 60
<< via1 >>
rect 804 2444 856 2496
rect 1844 2444 1896 2496
rect 44 2364 96 2416
rect 564 2364 616 2416
rect 1064 2364 1116 2416
rect 1584 2364 1636 2416
rect 2104 2364 2156 2416
rect 304 2304 356 2356
rect 1324 2304 1376 2356
rect 804 2064 856 2116
rect 1844 2064 1896 2116
rect 44 2004 96 2056
rect 564 2004 616 2056
rect 1064 2004 1116 2056
rect 1584 2004 1636 2056
rect 304 1924 356 1976
rect 1324 1924 1376 1976
rect 2104 2004 2156 2056
rect 804 1704 856 1756
rect 1844 1704 1896 1756
rect 44 1644 96 1696
rect 564 1644 616 1696
rect 1064 1644 1116 1696
rect 1584 1644 1636 1696
rect 304 1564 356 1616
rect 1324 1564 1376 1616
rect 2104 1644 2156 1696
rect 824 1344 876 1396
rect 1844 1344 1896 1396
rect 44 1284 96 1336
rect 564 1284 616 1336
rect 1064 1284 1116 1336
rect 1584 1284 1636 1336
rect 304 1204 356 1256
rect 1344 1204 1396 1256
rect 2104 1284 2156 1336
rect 804 984 856 1036
rect 1844 984 1896 1036
rect 44 904 96 956
rect 564 904 616 956
rect 1064 904 1116 956
rect 1584 904 1636 956
rect 304 844 356 896
rect 1324 844 1376 896
rect 2104 904 2156 956
rect 804 604 856 656
rect 1844 604 1896 656
rect 44 544 96 596
rect 564 544 616 596
rect 1064 544 1116 596
rect 1584 544 1636 596
rect 304 464 356 516
rect 1324 464 1376 516
rect 2104 544 2156 596
rect 804 244 856 296
rect 1844 244 1896 296
rect 44 184 96 236
rect 564 184 616 236
rect 1064 184 1116 236
rect 1584 184 1636 236
rect 304 104 356 156
rect 1324 104 1376 156
rect 2104 184 2156 236
<< metal2 >>
rect 800 2496 2320 2520
rect 800 2444 804 2496
rect 856 2480 1844 2496
rect 856 2444 860 2480
rect 800 2430 860 2444
rect 1840 2444 1844 2480
rect 1896 2480 2320 2496
rect 1896 2444 1900 2480
rect 1840 2430 1900 2444
rect 40 2418 100 2430
rect 40 2362 42 2418
rect 98 2362 100 2418
rect 560 2418 620 2430
rect 40 2350 100 2362
rect 300 2356 360 2370
rect 300 2320 304 2356
rect -120 2304 304 2320
rect 356 2320 360 2356
rect 560 2362 562 2418
rect 618 2362 620 2418
rect 560 2350 620 2362
rect 1060 2418 1120 2430
rect 1060 2362 1062 2418
rect 1118 2362 1120 2418
rect 1580 2418 1640 2430
rect 1060 2350 1120 2362
rect 1320 2356 1380 2370
rect 1320 2320 1324 2356
rect 356 2304 1324 2320
rect 1376 2304 1380 2356
rect 1580 2362 1582 2418
rect 1638 2362 1640 2418
rect 1580 2350 1640 2362
rect 2100 2418 2160 2430
rect 2100 2362 2102 2418
rect 2158 2362 2160 2418
rect 2100 2350 2160 2362
rect -120 2280 1380 2304
rect -120 2140 -40 2280
rect -120 2116 1900 2140
rect -120 2100 804 2116
rect -120 1580 -40 2100
rect 40 2058 100 2070
rect 40 2002 42 2058
rect 98 2002 100 2058
rect 40 1990 100 2002
rect 560 2058 620 2070
rect 560 2002 562 2058
rect 618 2002 620 2058
rect 800 2064 804 2100
rect 856 2100 1844 2116
rect 856 2064 860 2100
rect 800 2050 860 2064
rect 1060 2058 1120 2070
rect 560 1990 620 2002
rect 1060 2002 1062 2058
rect 1118 2002 1120 2058
rect 1060 1990 1120 2002
rect 1580 2058 1640 2070
rect 1580 2002 1582 2058
rect 1638 2002 1640 2058
rect 1840 2064 1844 2100
rect 1896 2064 1900 2116
rect 1840 2050 1900 2064
rect 2100 2058 2160 2070
rect 1580 1990 1640 2002
rect 2100 2002 2102 2058
rect 2158 2002 2160 2058
rect 2100 1990 2160 2002
rect 300 1976 360 1990
rect 300 1924 304 1976
rect 356 1940 360 1976
rect 1320 1976 1380 1990
rect 1320 1940 1324 1976
rect 356 1924 1324 1940
rect 1376 1940 1380 1976
rect 2240 1940 2320 2480
rect 1376 1924 2320 1940
rect 300 1900 2320 1924
rect 2240 1780 2320 1900
rect 800 1756 2320 1780
rect 40 1698 100 1710
rect 40 1642 42 1698
rect 98 1642 100 1698
rect 40 1630 100 1642
rect 560 1698 620 1710
rect 560 1642 562 1698
rect 618 1642 620 1698
rect 800 1704 804 1756
rect 856 1740 1844 1756
rect 856 1704 860 1740
rect 800 1690 860 1704
rect 1060 1698 1120 1710
rect 560 1630 620 1642
rect 1060 1642 1062 1698
rect 1118 1642 1120 1698
rect 1060 1630 1120 1642
rect 1580 1698 1640 1710
rect 1580 1642 1582 1698
rect 1638 1642 1640 1698
rect 1840 1704 1844 1740
rect 1896 1740 2320 1756
rect 1896 1704 1900 1740
rect 1840 1690 1900 1704
rect 2100 1698 2160 1710
rect 1580 1630 1640 1642
rect 2100 1642 2102 1698
rect 2158 1642 2160 1698
rect 2100 1630 2160 1642
rect 300 1616 360 1630
rect 300 1580 304 1616
rect -120 1564 304 1580
rect 356 1580 360 1616
rect 1320 1616 1380 1630
rect 1320 1580 1324 1616
rect 356 1564 1324 1580
rect 1376 1564 1380 1616
rect -120 1540 1380 1564
rect -120 1420 -40 1540
rect -120 1396 1900 1420
rect -120 1380 824 1396
rect -120 860 -40 1380
rect 40 1338 100 1350
rect 40 1282 42 1338
rect 98 1282 100 1338
rect 40 1270 100 1282
rect 560 1338 620 1350
rect 560 1282 562 1338
rect 618 1282 620 1338
rect 820 1344 824 1380
rect 876 1380 1844 1396
rect 876 1344 880 1380
rect 820 1330 880 1344
rect 1060 1338 1120 1350
rect 560 1270 620 1282
rect 1060 1282 1062 1338
rect 1118 1282 1120 1338
rect 1060 1270 1120 1282
rect 1580 1338 1640 1350
rect 1580 1282 1582 1338
rect 1638 1282 1640 1338
rect 1840 1344 1844 1380
rect 1896 1344 1900 1396
rect 1840 1330 1900 1344
rect 2100 1338 2160 1350
rect 1580 1270 1640 1282
rect 2100 1282 2102 1338
rect 2158 1282 2160 1338
rect 2100 1270 2160 1282
rect 300 1256 360 1270
rect 300 1204 304 1256
rect 356 1220 360 1256
rect 1340 1256 1400 1270
rect 1340 1220 1344 1256
rect 356 1204 1344 1220
rect 1396 1220 1400 1256
rect 2240 1220 2320 1740
rect 1396 1204 2320 1220
rect 300 1180 2320 1204
rect 2240 1060 2320 1180
rect 800 1036 2320 1060
rect 800 984 804 1036
rect 856 1020 1844 1036
rect 856 984 860 1020
rect 800 970 860 984
rect 1840 984 1844 1020
rect 1896 1020 2320 1036
rect 1896 984 1900 1020
rect 1840 970 1900 984
rect 40 958 100 970
rect 40 902 42 958
rect 98 902 100 958
rect 560 958 620 970
rect 40 890 100 902
rect 300 896 360 910
rect 300 860 304 896
rect -120 844 304 860
rect 356 860 360 896
rect 560 902 562 958
rect 618 902 620 958
rect 560 890 620 902
rect 1060 958 1120 970
rect 1060 902 1062 958
rect 1118 902 1120 958
rect 1580 958 1640 970
rect 1060 890 1120 902
rect 1320 896 1380 910
rect 1320 860 1324 896
rect 356 844 1324 860
rect 1376 844 1380 896
rect 1580 902 1582 958
rect 1638 902 1640 958
rect 1580 890 1640 902
rect 2100 958 2160 970
rect 2100 902 2102 958
rect 2158 902 2160 958
rect 2100 890 2160 902
rect -120 820 1380 844
rect -120 680 -40 820
rect -120 656 1900 680
rect -120 640 804 656
rect -120 120 -40 640
rect 40 598 100 610
rect 40 542 42 598
rect 98 542 100 598
rect 40 530 100 542
rect 560 598 620 610
rect 560 542 562 598
rect 618 542 620 598
rect 800 604 804 640
rect 856 640 1844 656
rect 856 604 860 640
rect 800 590 860 604
rect 1060 598 1120 610
rect 560 530 620 542
rect 1060 542 1062 598
rect 1118 542 1120 598
rect 1060 530 1120 542
rect 1580 598 1640 610
rect 1580 542 1582 598
rect 1638 542 1640 598
rect 1840 604 1844 640
rect 1896 604 1900 656
rect 1840 590 1900 604
rect 2100 598 2160 610
rect 1580 530 1640 542
rect 2100 542 2102 598
rect 2158 542 2160 598
rect 2100 530 2160 542
rect 300 516 360 530
rect 300 464 304 516
rect 356 480 360 516
rect 1320 516 1380 530
rect 1320 480 1324 516
rect 356 464 1324 480
rect 1376 480 1380 516
rect 2240 480 2320 1020
rect 1376 464 2320 480
rect 300 440 2320 464
rect 2240 320 2320 440
rect 800 296 2320 320
rect 40 238 100 250
rect 40 182 42 238
rect 98 182 100 238
rect 40 170 100 182
rect 560 238 620 250
rect 560 182 562 238
rect 618 182 620 238
rect 800 244 804 296
rect 856 280 1844 296
rect 856 244 860 280
rect 800 230 860 244
rect 1060 238 1120 250
rect 560 170 620 182
rect 1060 182 1062 238
rect 1118 182 1120 238
rect 1060 170 1120 182
rect 1580 238 1640 250
rect 1580 182 1582 238
rect 1638 182 1640 238
rect 1840 244 1844 280
rect 1896 280 2320 296
rect 1896 244 1900 280
rect 1840 230 1900 244
rect 2100 238 2160 250
rect 1580 170 1640 182
rect 2100 182 2102 238
rect 2158 182 2160 238
rect 2100 170 2160 182
rect 300 156 360 170
rect 300 120 304 156
rect -120 104 304 120
rect 356 120 360 156
rect 1320 156 1380 170
rect 1320 120 1324 156
rect 356 104 1324 120
rect 1376 104 1380 156
rect -120 80 1380 104
<< via2 >>
rect 42 2416 98 2418
rect 42 2364 44 2416
rect 44 2364 96 2416
rect 96 2364 98 2416
rect 42 2362 98 2364
rect 562 2416 618 2418
rect 562 2364 564 2416
rect 564 2364 616 2416
rect 616 2364 618 2416
rect 562 2362 618 2364
rect 1062 2416 1118 2418
rect 1062 2364 1064 2416
rect 1064 2364 1116 2416
rect 1116 2364 1118 2416
rect 1062 2362 1118 2364
rect 1582 2416 1638 2418
rect 1582 2364 1584 2416
rect 1584 2364 1636 2416
rect 1636 2364 1638 2416
rect 1582 2362 1638 2364
rect 2102 2416 2158 2418
rect 2102 2364 2104 2416
rect 2104 2364 2156 2416
rect 2156 2364 2158 2416
rect 2102 2362 2158 2364
rect 42 2056 98 2058
rect 42 2004 44 2056
rect 44 2004 96 2056
rect 96 2004 98 2056
rect 42 2002 98 2004
rect 562 2056 618 2058
rect 562 2004 564 2056
rect 564 2004 616 2056
rect 616 2004 618 2056
rect 562 2002 618 2004
rect 1062 2056 1118 2058
rect 1062 2004 1064 2056
rect 1064 2004 1116 2056
rect 1116 2004 1118 2056
rect 1062 2002 1118 2004
rect 1582 2056 1638 2058
rect 1582 2004 1584 2056
rect 1584 2004 1636 2056
rect 1636 2004 1638 2056
rect 1582 2002 1638 2004
rect 2102 2056 2158 2058
rect 2102 2004 2104 2056
rect 2104 2004 2156 2056
rect 2156 2004 2158 2056
rect 2102 2002 2158 2004
rect 42 1696 98 1698
rect 42 1644 44 1696
rect 44 1644 96 1696
rect 96 1644 98 1696
rect 42 1642 98 1644
rect 562 1696 618 1698
rect 562 1644 564 1696
rect 564 1644 616 1696
rect 616 1644 618 1696
rect 562 1642 618 1644
rect 1062 1696 1118 1698
rect 1062 1644 1064 1696
rect 1064 1644 1116 1696
rect 1116 1644 1118 1696
rect 1062 1642 1118 1644
rect 1582 1696 1638 1698
rect 1582 1644 1584 1696
rect 1584 1644 1636 1696
rect 1636 1644 1638 1696
rect 1582 1642 1638 1644
rect 2102 1696 2158 1698
rect 2102 1644 2104 1696
rect 2104 1644 2156 1696
rect 2156 1644 2158 1696
rect 2102 1642 2158 1644
rect 42 1336 98 1338
rect 42 1284 44 1336
rect 44 1284 96 1336
rect 96 1284 98 1336
rect 42 1282 98 1284
rect 562 1336 618 1338
rect 562 1284 564 1336
rect 564 1284 616 1336
rect 616 1284 618 1336
rect 562 1282 618 1284
rect 1062 1336 1118 1338
rect 1062 1284 1064 1336
rect 1064 1284 1116 1336
rect 1116 1284 1118 1336
rect 1062 1282 1118 1284
rect 1582 1336 1638 1338
rect 1582 1284 1584 1336
rect 1584 1284 1636 1336
rect 1636 1284 1638 1336
rect 1582 1282 1638 1284
rect 2102 1336 2158 1338
rect 2102 1284 2104 1336
rect 2104 1284 2156 1336
rect 2156 1284 2158 1336
rect 2102 1282 2158 1284
rect 42 956 98 958
rect 42 904 44 956
rect 44 904 96 956
rect 96 904 98 956
rect 42 902 98 904
rect 562 956 618 958
rect 562 904 564 956
rect 564 904 616 956
rect 616 904 618 956
rect 562 902 618 904
rect 1062 956 1118 958
rect 1062 904 1064 956
rect 1064 904 1116 956
rect 1116 904 1118 956
rect 1062 902 1118 904
rect 1582 956 1638 958
rect 1582 904 1584 956
rect 1584 904 1636 956
rect 1636 904 1638 956
rect 1582 902 1638 904
rect 2102 956 2158 958
rect 2102 904 2104 956
rect 2104 904 2156 956
rect 2156 904 2158 956
rect 2102 902 2158 904
rect 42 596 98 598
rect 42 544 44 596
rect 44 544 96 596
rect 96 544 98 596
rect 42 542 98 544
rect 562 596 618 598
rect 562 544 564 596
rect 564 544 616 596
rect 616 544 618 596
rect 562 542 618 544
rect 1062 596 1118 598
rect 1062 544 1064 596
rect 1064 544 1116 596
rect 1116 544 1118 596
rect 1062 542 1118 544
rect 1582 596 1638 598
rect 1582 544 1584 596
rect 1584 544 1636 596
rect 1636 544 1638 596
rect 1582 542 1638 544
rect 2102 596 2158 598
rect 2102 544 2104 596
rect 2104 544 2156 596
rect 2156 544 2158 596
rect 2102 542 2158 544
rect 42 236 98 238
rect 42 184 44 236
rect 44 184 96 236
rect 96 184 98 236
rect 42 182 98 184
rect 562 236 618 238
rect 562 184 564 236
rect 564 184 616 236
rect 616 184 618 236
rect 562 182 618 184
rect 1062 236 1118 238
rect 1062 184 1064 236
rect 1064 184 1116 236
rect 1116 184 1118 236
rect 1062 182 1118 184
rect 1582 236 1638 238
rect 1582 184 1584 236
rect 1584 184 1636 236
rect 1636 184 1638 236
rect 1582 182 1638 184
rect 2102 236 2158 238
rect 2102 184 2104 236
rect 2104 184 2156 236
rect 2156 184 2158 236
rect 2102 182 2158 184
<< metal3 >>
rect 40 2425 100 2500
rect 560 2425 620 2500
rect 1060 2425 1120 2500
rect 1580 2425 1640 2500
rect 2100 2425 2160 2500
rect 30 2418 110 2425
rect 30 2362 42 2418
rect 98 2362 110 2418
rect 30 2355 110 2362
rect 550 2418 630 2425
rect 550 2362 562 2418
rect 618 2362 630 2418
rect 550 2355 630 2362
rect 1050 2418 1130 2425
rect 1050 2362 1062 2418
rect 1118 2362 1130 2418
rect 1050 2355 1130 2362
rect 1570 2418 1650 2425
rect 1570 2362 1582 2418
rect 1638 2362 1650 2418
rect 1570 2355 1650 2362
rect 2090 2418 2170 2425
rect 2090 2362 2102 2418
rect 2158 2362 2170 2418
rect 2090 2355 2170 2362
rect 40 2065 100 2355
rect 560 2065 620 2355
rect 1060 2065 1120 2355
rect 1580 2065 1640 2355
rect 2100 2065 2160 2355
rect 30 2058 110 2065
rect 30 2002 42 2058
rect 98 2002 110 2058
rect 30 1995 110 2002
rect 550 2058 630 2065
rect 550 2002 562 2058
rect 618 2002 630 2058
rect 550 1995 630 2002
rect 1050 2058 1130 2065
rect 1050 2002 1062 2058
rect 1118 2002 1130 2058
rect 1050 1995 1130 2002
rect 1570 2058 1650 2065
rect 1570 2002 1582 2058
rect 1638 2002 1650 2058
rect 1570 1995 1650 2002
rect 2090 2058 2170 2065
rect 2090 2002 2102 2058
rect 2158 2002 2170 2058
rect 2090 1995 2170 2002
rect 40 1705 100 1995
rect 560 1705 620 1995
rect 1060 1705 1120 1995
rect 1580 1705 1640 1995
rect 2100 1705 2160 1995
rect 30 1698 110 1705
rect 30 1642 42 1698
rect 98 1642 110 1698
rect 30 1635 110 1642
rect 550 1698 630 1705
rect 550 1642 562 1698
rect 618 1642 630 1698
rect 550 1635 630 1642
rect 1050 1698 1130 1705
rect 1050 1642 1062 1698
rect 1118 1642 1130 1698
rect 1050 1635 1130 1642
rect 1570 1698 1650 1705
rect 1570 1642 1582 1698
rect 1638 1642 1650 1698
rect 1570 1635 1650 1642
rect 2090 1698 2170 1705
rect 2090 1642 2102 1698
rect 2158 1642 2170 1698
rect 2090 1635 2170 1642
rect 40 1345 100 1635
rect 560 1345 620 1635
rect 1060 1345 1120 1635
rect 1580 1345 1640 1635
rect 2100 1345 2160 1635
rect 30 1340 110 1345
rect 550 1340 630 1345
rect 1050 1340 1130 1345
rect 1570 1340 1650 1345
rect 2090 1340 2170 1345
rect -120 1338 2320 1340
rect -120 1282 42 1338
rect 98 1282 562 1338
rect 618 1282 1062 1338
rect 1118 1282 1582 1338
rect 1638 1282 2102 1338
rect 2158 1282 2320 1338
rect -120 1280 2320 1282
rect 30 1275 110 1280
rect 550 1275 630 1280
rect 1050 1275 1130 1280
rect 1570 1275 1650 1280
rect 2090 1275 2170 1280
rect 40 965 100 1275
rect 560 965 620 1275
rect 1060 965 1120 1275
rect 1580 965 1640 1275
rect 2100 965 2160 1275
rect 30 958 110 965
rect 30 902 42 958
rect 98 902 110 958
rect 30 895 110 902
rect 550 958 630 965
rect 550 902 562 958
rect 618 902 630 958
rect 550 895 630 902
rect 1050 958 1130 965
rect 1050 902 1062 958
rect 1118 902 1130 958
rect 1050 895 1130 902
rect 1570 958 1650 965
rect 1570 902 1582 958
rect 1638 902 1650 958
rect 1570 895 1650 902
rect 2090 958 2170 965
rect 2090 902 2102 958
rect 2158 902 2170 958
rect 2090 895 2170 902
rect 40 605 100 895
rect 560 605 620 895
rect 1060 605 1120 895
rect 1580 605 1640 895
rect 2100 605 2160 895
rect 30 598 110 605
rect 30 542 42 598
rect 98 542 110 598
rect 30 535 110 542
rect 550 598 630 605
rect 550 542 562 598
rect 618 542 630 598
rect 550 535 630 542
rect 1050 598 1130 605
rect 1050 542 1062 598
rect 1118 542 1130 598
rect 1050 535 1130 542
rect 1570 598 1650 605
rect 1570 542 1582 598
rect 1638 542 1650 598
rect 1570 535 1650 542
rect 2090 598 2170 605
rect 2090 542 2102 598
rect 2158 542 2170 598
rect 2090 535 2170 542
rect 40 245 100 535
rect 560 245 620 535
rect 1060 245 1120 535
rect 1580 245 1640 535
rect 2100 245 2160 535
rect 30 238 110 245
rect 30 182 42 238
rect 98 182 110 238
rect 30 175 110 182
rect 550 238 630 245
rect 550 182 562 238
rect 618 182 630 238
rect 550 175 630 182
rect 1050 238 1130 245
rect 1050 182 1062 238
rect 1118 182 1130 238
rect 1050 175 1130 182
rect 1570 238 1650 245
rect 1570 182 1582 238
rect 1638 182 1650 238
rect 1570 175 1650 182
rect 2090 238 2170 245
rect 2090 182 2102 238
rect 2158 182 2170 238
rect 2090 175 2170 182
rect 40 100 100 175
rect 560 100 620 175
rect 1060 100 1120 175
rect 1580 100 1640 175
rect 2100 100 2160 175
use sky130_fd_pr__pfet_01v8_lvt_8URDWJ  sky130_fd_pr__pfet_01v8_lvt_8URDWJ_0
timestamp 1663011646
transform 1 0 1097 0 1 1260
box -1097 -1260 1097 1292
<< labels >>
flabel nwell s 300 2540 360 2620 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1340 2540 1400 2620 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 820 2160 880 2240 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1840 2140 1900 2220 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 280 1780 340 1860 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1340 1800 1400 1880 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 820 1400 880 1480 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1840 1400 1900 1480 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 300 1040 360 1120 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1340 1060 1400 1140 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 780 680 840 760 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1860 680 1920 760 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 280 300 340 380 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 1320 300 1380 380 0 FreeSans 1000 0 0 0 A
port 1 nsew
flabel nwell s 820 2520 880 2600 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1840 2520 1900 2600 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 300 2140 360 2220 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1340 2140 1400 2220 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 820 1780 880 1860 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1860 1780 1920 1860 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 280 1400 340 1480 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1340 1420 1400 1500 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 820 1060 880 1140 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1840 1060 1900 1140 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 300 700 360 780 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1340 680 1400 760 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 820 320 880 400 0 FreeSans 1000 0 0 0 B
port 2 nsew
flabel nwell s 1840 320 1900 400 0 FreeSans 1000 0 0 0 B
port 2 nsew
<< end >>
