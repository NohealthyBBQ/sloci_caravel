magic
tech sky130A
magscale 1 2
timestamp 1669931957
<< metal1 >>
rect 14920 682870 15420 682910
rect 14920 682040 14960 682870
rect 15390 682040 15420 682870
rect 14920 668280 15420 682040
rect 14920 668180 23410 668280
rect 14920 668100 23840 668180
rect 14920 668060 23410 668100
rect 14920 433640 15420 668060
rect 55960 662600 56100 662620
rect 55960 662500 55980 662600
rect 56080 662500 56100 662600
rect 55960 662480 56100 662500
rect 56200 661680 56340 661700
rect 56200 661580 56220 661680
rect 56320 661580 56340 661680
rect 56200 661560 56340 661580
rect 56480 661080 56620 661100
rect 56480 660980 56500 661080
rect 56600 660980 56620 661080
rect 56480 660960 56620 660980
rect 56720 660560 56860 660580
rect 56720 660460 56740 660560
rect 56840 660460 56860 660560
rect 56720 660440 56860 660460
rect 56980 660200 57120 660220
rect 56980 660100 57000 660200
rect 57100 660100 57120 660200
rect 56980 660080 57120 660100
rect 14920 433480 144980 433640
rect 144900 432740 144980 433480
rect 55960 400380 58040 400400
rect 55960 400300 55980 400380
rect 56080 400300 57920 400380
rect 58020 400300 58040 400380
rect 55960 400280 58040 400300
rect 139220 400380 139340 400400
rect 139220 400300 139240 400380
rect 139220 400280 139340 400300
rect 56200 400120 58040 400140
rect 56200 400040 56220 400120
rect 56320 400040 57920 400120
rect 58020 400040 58040 400120
rect 56200 400020 58040 400040
rect 138320 400120 138460 400140
rect 138320 400040 138340 400120
rect 138440 400040 138460 400120
rect 138320 400020 138460 400040
rect 56480 399860 58040 399880
rect 56480 399780 56500 399860
rect 56600 399780 57920 399860
rect 58020 399780 58040 399860
rect 56480 399760 58040 399780
rect 137720 399860 137860 399880
rect 137720 399780 137740 399860
rect 137840 399780 137860 399860
rect 137720 399760 137860 399780
rect 56720 399600 58040 399620
rect 56720 399520 56740 399600
rect 56840 399520 57920 399600
rect 58020 399520 58040 399600
rect 56720 399500 58040 399520
rect 137180 399600 137320 399620
rect 137180 399520 137200 399600
rect 137300 399520 137320 399600
rect 137180 399500 137320 399520
rect 136820 399340 136960 399360
rect 136820 399260 136840 399340
rect 136940 399260 136960 399340
rect 136820 399240 136960 399260
<< via1 >>
rect 14960 682040 15390 682870
rect 55980 662500 56080 662600
rect 56220 661580 56320 661680
rect 56500 660980 56600 661080
rect 56740 660460 56840 660560
rect 57000 660100 57100 660200
rect 55980 400300 56080 400380
rect 57920 400300 58020 400380
rect 139240 400300 139340 400380
rect 56220 400040 56320 400120
rect 57920 400040 58020 400120
rect 138340 400040 138440 400120
rect 56500 399780 56600 399860
rect 57920 399780 58020 399860
rect 137740 399780 137840 399860
rect 56740 399520 56840 399600
rect 57920 399520 58020 399600
rect 137200 399520 137300 399600
rect 136840 399260 136940 399340
<< metal2 >>
rect 14920 682870 15420 682910
rect 14920 682040 14960 682870
rect 15390 682040 15420 682870
rect 14920 681990 15420 682040
rect 23190 671610 25400 671620
rect 23190 671440 23210 671610
rect 23370 671440 25400 671610
rect 23190 671420 25400 671440
rect 55960 662600 56100 662700
rect 55960 662500 55980 662600
rect 56080 662500 56100 662600
rect 55960 400380 56100 662500
rect 55960 400300 55980 400380
rect 56080 400300 56100 400380
rect 55960 292200 56100 400300
rect 56200 661680 56340 661700
rect 56200 661580 56220 661680
rect 56320 661580 56340 661680
rect 56200 400120 56340 661580
rect 56200 400040 56220 400120
rect 56320 400040 56340 400120
rect 56200 335220 56340 400040
rect 56480 661080 56620 661100
rect 56480 660980 56500 661080
rect 56600 660980 56620 661080
rect 56480 399860 56620 660980
rect 56480 399780 56500 399860
rect 56600 399780 56620 399860
rect 56480 378460 56620 399780
rect 56720 660560 56860 660580
rect 56720 660460 56740 660560
rect 56840 660460 56860 660560
rect 56720 421660 56860 660460
rect 56720 421520 56740 421660
rect 56840 421520 56860 421660
rect 56720 399600 56860 421520
rect 56720 399520 56740 399600
rect 56840 399520 56860 399600
rect 56720 399500 56860 399520
rect 56980 660200 57120 660220
rect 56980 660100 57000 660200
rect 57100 660100 57120 660200
rect 56980 466080 57120 660100
rect 238000 591000 246800 592200
rect 238000 582000 239000 591000
rect 246000 582000 246800 591000
rect 238000 580200 246800 582000
rect 246300 579400 246700 580200
rect 56980 465940 57000 466080
rect 57100 465940 57120 466080
rect 56980 399360 57120 465940
rect 148000 435600 149000 436000
rect 148000 434400 148200 435600
rect 148800 434400 149000 435600
rect 148000 434000 149000 434400
rect 148200 430920 148420 434000
rect 57900 400380 139360 400400
rect 57900 400300 57920 400380
rect 58020 400300 139240 400380
rect 139340 400300 139360 400380
rect 57900 400280 139360 400300
rect 57900 400120 138460 400140
rect 57900 400040 57920 400120
rect 58020 400040 138340 400120
rect 138440 400040 138460 400120
rect 57900 400020 138460 400040
rect 57900 399860 137860 399880
rect 57900 399780 57920 399860
rect 58020 399780 137740 399860
rect 137840 399780 137860 399860
rect 57900 399760 137860 399780
rect 57900 399600 137320 399620
rect 57900 399520 57920 399600
rect 58020 399520 137200 399600
rect 137300 399520 137320 399600
rect 57900 399500 137320 399520
rect 56980 399340 136960 399360
rect 56980 399260 136840 399340
rect 136940 399260 136960 399340
rect 56980 399240 136960 399260
rect 56480 378320 56500 378460
rect 56600 378320 56620 378460
rect 56480 378300 56620 378320
rect 56200 335080 56220 335220
rect 56320 335080 56340 335220
rect 56200 335060 56340 335080
rect 55960 291860 55980 292000
rect 56080 291860 56100 292000
rect 55960 291840 56100 291860
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 14960 682040 15390 682870
rect 23210 671440 23370 671610
rect 56740 421520 56840 421660
rect 239000 582000 246000 591000
rect 57000 465940 57100 466080
rect 148200 434400 148800 435600
rect 56500 378320 56600 378460
rect 56220 335080 56320 335220
rect 55980 291860 56080 292000
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 704000 125194 704800
rect 17070 689360 19380 702300
rect 68470 689480 70760 702300
rect 42500 689440 70760 689480
rect 17070 689330 26050 689360
rect 17070 688210 41870 689330
rect 42500 688410 42560 689440
rect 43180 688410 70760 689440
rect 42500 688360 70760 688410
rect 17070 688200 26050 688210
rect -800 682910 1700 685242
rect -800 682870 15420 682910
rect -800 682040 14960 682870
rect 15390 682040 15420 682870
rect -800 681990 15420 682040
rect -800 680242 1700 681990
rect 40710 680350 41870 688210
rect 40720 679110 41870 680350
rect 40720 677240 41720 677320
rect 40720 676130 40770 677240
rect 41640 676130 41720 677240
rect 40720 676080 41720 676130
rect 23190 671610 23390 671620
rect 23190 671440 23210 671610
rect 23370 671440 23390 671610
rect 23190 669080 23390 671440
rect 23190 668680 23210 669080
rect 23370 668680 23390 669080
rect 23190 668640 23390 668680
rect 310 648642 1780 648730
rect -800 648600 1780 648642
rect -800 648200 5000 648600
rect -800 643842 2200 648200
rect 246 638642 2200 643842
rect -800 634200 2200 638642
rect 4600 634200 5000 648200
rect -800 633842 5000 634200
rect 246 633838 5000 633842
rect 1800 633800 5000 633838
rect 120000 606000 126000 704000
rect 165594 702300 170594 704800
rect 170894 702300 173094 704800
rect 173394 703000 175594 704800
rect 173394 702300 175600 703000
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 222594 702300 224794 704800
rect 225094 702300 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 324294 702300 326494 704800
rect 326794 702300 328994 704800
rect 329294 702300 334294 704800
rect 413394 702412 418394 704800
rect 173400 702200 175600 702300
rect 413334 702000 413344 702412
rect 418488 702000 418498 702412
rect 465394 702376 470394 704800
rect 465328 700564 471268 702376
rect 510594 702340 515394 704800
rect 520594 702340 525394 704800
rect 566594 702300 571594 704800
rect 582300 677984 584800 682984
rect 582296 644584 583800 644600
rect 582296 639784 584800 644584
rect 582296 634584 583800 639784
rect 582296 629800 584800 634584
rect 582340 629784 584800 629800
rect 288200 606000 289800 606600
rect 21990 605800 24010 606000
rect 21990 605000 22400 605800
rect 23600 605000 24010 605800
rect 21990 604000 24010 605000
rect 120000 604000 290000 606000
rect 22000 602000 24000 604000
rect 22000 600000 287600 602000
rect 147000 595800 285400 596000
rect 147000 594200 148200 595800
rect 148800 594200 285400 595800
rect 147000 594000 285400 594200
rect 238990 591000 246010 591005
rect 164000 590000 239000 591000
rect 164000 583000 165000 590000
rect 182000 583000 239000 590000
rect 164000 582000 239000 583000
rect 246000 582000 246010 591000
rect 238990 581995 246010 582000
rect 85400 580000 245900 581400
rect 283800 580600 285400 594000
rect 286000 580600 287600 600000
rect 288200 580600 289800 604000
rect 290506 594136 292488 595526
rect 290546 580594 292130 594136
rect 293590 592863 295448 592882
rect 292774 591450 295448 592863
rect 292774 580566 294378 591450
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 581366 587220 583814 587614
rect 581366 587108 584800 587220
rect 581366 587056 583814 587108
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 564220 1660 564242
rect -800 564080 4430 564220
rect -800 559570 860 564080
rect 4260 559570 4430 564080
rect -800 559442 4430 559570
rect 680 555000 4430 559442
rect 680 554242 1000 555000
rect -800 550000 1000 554242
rect 4000 550000 4430 555000
rect -800 549442 4430 550000
rect 680 549410 4430 549442
rect 85400 511800 86800 580000
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 400 511642 86800 511800
rect -800 511530 86800 511642
rect 400 511200 86800 511530
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 583520 495322 584800 495434
rect 583520 494140 584800 494252
rect -800 468308 480 468420
rect 163400 467800 200000 468000
rect -800 467126 480 467238
rect 163400 466200 198200 467800
rect 199800 466200 200000 467800
rect 280 466080 57120 466100
rect 280 466056 57000 466080
rect -800 465944 57000 466056
rect 280 465940 57000 465944
rect 57100 465940 57120 466080
rect 280 465920 57120 465940
rect 163400 466000 200000 466200
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 148000 435800 149000 436000
rect 148000 434200 148200 435800
rect 148800 434200 149000 435800
rect 148000 434000 149000 434200
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect 360 421660 56860 421680
rect 360 421652 56740 421660
rect -800 421540 56740 421652
rect 360 421520 56740 421540
rect 56840 421520 56860 421660
rect 360 421500 56860 421520
rect -800 420358 480 420470
rect -800 419176 480 419288
rect 163400 415700 164900 466000
rect 583520 455628 584800 455740
rect 583520 454446 584800 454558
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 583520 449718 584800 449830
rect 152900 415200 154200 415700
rect 155900 415200 164900 415700
rect 152900 414870 153400 415200
rect 152900 414440 152960 414870
rect 153360 414440 153400 414870
rect 152900 414400 153400 414440
rect 158890 414870 164900 414900
rect 158890 414440 158950 414870
rect 159350 414440 164900 414870
rect 158890 414400 164900 414440
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect 400 378460 56620 378480
rect 400 378430 56500 378460
rect -800 378320 56500 378430
rect 56600 378320 56620 378460
rect -800 378318 56620 378320
rect 400 378300 56620 378318
rect -800 377136 480 377248
rect -800 375954 480 376066
rect 163400 362000 164900 414400
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 163400 361800 200000 362000
rect 163400 360200 198200 361800
rect 199800 360200 200000 361800
rect 583520 361238 584800 361350
rect 163400 360000 200000 360200
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect 260 335220 56340 335240
rect 260 335208 56220 335220
rect -800 335096 56220 335208
rect 260 335080 56220 335096
rect 56320 335080 56340 335220
rect 260 335060 56340 335080
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect 200 295532 800 295600
rect -800 295420 800 295532
rect 200 295400 800 295420
rect 200 294350 800 294400
rect -800 294238 800 294350
rect 200 294200 800 294238
rect -800 293056 480 293168
rect 400 292000 56100 292020
rect 400 291986 55980 292000
rect -800 291874 55980 291986
rect 400 291860 55980 291874
rect 56080 291860 56100 292000
rect 400 291840 56100 291860
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect 4160 219700 17580 219880
rect 1660 219688 17580 219700
rect -800 219500 17580 219688
rect -800 214888 11340 219500
rect 1660 210740 11340 214888
rect 17140 210740 17580 219500
rect 1660 210380 17580 210740
rect 1660 209688 5520 210380
rect -800 204900 5520 209688
rect -800 204888 1660 204900
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect 982 177688 1680 177690
rect -800 172888 1680 177688
rect 982 172880 1680 172888
rect -800 167680 1660 167688
rect -800 162890 1680 167680
rect -800 162888 1660 162890
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 42560 688410 43180 689440
rect 40770 676130 41640 677240
rect 23210 668680 23370 669080
rect 2200 634200 4600 648200
rect 413344 702000 418488 702412
rect 22400 605000 23600 605800
rect 148200 594200 148800 595800
rect 165000 583000 182000 590000
rect 860 559570 4260 564080
rect 1000 550000 4000 555000
rect 198200 466200 199800 467800
rect 148200 435600 148800 435800
rect 148200 434400 148800 435600
rect 148200 434200 148800 434400
rect 152960 414440 153360 414870
rect 158950 414440 159350 414870
rect 198200 360200 199800 361800
rect 11340 210740 17140 219500
<< metal4 >>
rect 165594 703000 170594 704800
rect 175894 703000 180894 704800
rect 42500 689440 43450 689470
rect 42500 688410 42560 689440
rect 43180 688410 43450 689440
rect 42500 677320 43450 688410
rect 40720 677240 43450 677320
rect 40720 676130 40770 677240
rect 41640 676130 43450 677240
rect 40720 676090 43450 676130
rect 40720 676080 43220 676090
rect 60220 676010 65450 676030
rect 56870 675370 65450 676010
rect 23190 669080 23390 669110
rect 23190 668680 23210 669080
rect 23370 668680 23390 669080
rect 1800 648200 5000 648600
rect 1800 634200 2200 648200
rect 4600 634200 5000 648200
rect 1800 633800 5000 634200
rect 23190 619600 23390 668680
rect 25400 662640 27800 663400
rect 25400 633690 28120 662640
rect 32000 658600 39600 659000
rect 32000 656800 32200 658600
rect 39200 656800 39600 658600
rect 25400 631490 28200 633690
rect 22600 611800 23400 619600
rect 22200 605800 23800 611800
rect 22200 605000 22400 605800
rect 23600 605000 23800 605800
rect 22200 604800 23800 605000
rect 690 564080 4450 564270
rect 690 559570 860 564080
rect 4260 559570 4450 564080
rect 690 559400 4450 559570
rect 25400 564000 28000 631490
rect 32000 620900 39600 656800
rect 32000 618600 39650 620900
rect 32100 613600 39650 618600
rect 999 555000 4001 555001
rect 999 550000 1000 555000
rect 4000 550000 4001 555000
rect 25400 550600 25800 564000
rect 27600 550600 28000 564000
rect 25400 550200 28000 550600
rect 999 549999 4001 550000
rect 30150 418600 39650 613600
rect 60600 564000 65400 675370
rect 165000 664570 182000 703000
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 413343 702412 418489 702413
rect 413343 702000 413344 702412
rect 418488 702000 418489 702412
rect 413343 701999 418489 702000
rect 165000 659662 168158 664570
rect 179872 659662 182000 664570
rect 148000 595800 149000 596000
rect 148000 594200 148200 595800
rect 148800 594200 149000 595800
rect 60600 550400 61000 564000
rect 65000 550400 65400 564000
rect 60600 550000 65400 550400
rect 126400 563600 131200 564000
rect 126400 550400 126800 563600
rect 130800 550400 131200 563600
rect 30150 409800 30600 418600
rect 39000 409800 39650 418600
rect 30150 219860 39650 409800
rect 126400 429800 131200 550400
rect 148000 435800 149000 594200
rect 165000 590001 182000 659662
rect 305500 645000 316500 646500
rect 164999 590000 182001 590001
rect 164999 583000 165000 590000
rect 182000 583000 182001 590000
rect 164999 582999 182001 583000
rect 238000 584000 248000 636000
rect 305500 637000 307000 645000
rect 315000 637000 316500 645000
rect 238000 580000 260000 584000
rect 305500 580300 316500 637000
rect 238200 570900 240100 574000
rect 258800 571400 260000 580000
rect 238200 568100 239300 570900
rect 238200 563700 240200 568100
rect 239700 558000 240200 563700
rect 263600 557900 316600 558100
rect 198000 467800 200000 468000
rect 198000 466200 198200 467800
rect 199800 466200 200000 467800
rect 198000 466000 200000 466200
rect 148000 434200 148200 435800
rect 148800 434200 149000 435800
rect 148000 434000 149000 434200
rect 126400 428200 139400 429800
rect 126400 399000 131200 428200
rect 152900 414870 159400 414900
rect 152900 414440 152960 414870
rect 153360 414440 158950 414870
rect 159350 414440 159400 414870
rect 152900 414400 159400 414440
rect 126400 397800 152800 399000
rect 198000 361800 200000 362000
rect 198000 360200 198200 361800
rect 199800 360200 200000 361800
rect 198000 360000 200000 360200
rect 10880 219500 39650 219860
rect 10880 210740 11340 219500
rect 17140 214040 39650 219500
rect 17140 210740 39640 214040
rect 10880 210360 39640 210740
<< via4 >>
rect 2200 635400 4600 646600
rect 32200 656800 39200 658600
rect 860 559570 4260 564080
rect 1000 550000 4000 555000
rect 25800 550600 27600 564000
rect 168158 659662 179872 664570
rect 61000 550400 65000 564000
rect 126800 550400 130800 563600
rect 30600 409800 39000 418600
rect 238000 636000 248000 644000
rect 307000 637000 315000 645000
rect 238200 558000 239700 563700
rect 263600 556400 316600 557900
rect 198200 466200 199800 467800
rect 198200 360200 199800 361800
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 329294 702300 334294 704800
rect 32000 659200 33600 675200
rect 35600 659200 36200 675200
rect 38800 659200 39400 675200
rect 42200 659200 43800 675200
rect 168134 664570 179896 664594
rect 45800 659200 46400 660800
rect 168134 659662 168158 664570
rect 179872 659662 179896 664570
rect 168134 659638 179896 659662
rect 32000 658600 46400 659200
rect 32000 656800 32200 658600
rect 39200 656800 46400 658600
rect 32000 656400 46400 656800
rect 72976 647000 79024 647024
rect 1800 646600 320000 647000
rect 1800 635400 2200 646600
rect 4600 645000 320000 646600
rect 4600 644000 307000 645000
rect 4600 636000 238000 644000
rect 248000 637000 307000 644000
rect 315000 637000 320000 645000
rect 248000 636000 320000 637000
rect 4600 635400 320000 636000
rect 1800 635000 320000 635400
rect 72976 634976 79024 635000
rect 60760 564330 65600 564340
rect 28810 564320 65600 564330
rect 1770 564270 65600 564320
rect 690 564080 65600 564270
rect 690 559570 860 564080
rect 4260 564000 65600 564080
rect 4260 559570 25800 564000
rect 690 559400 25800 559570
rect 1000 555024 25800 559400
rect 976 555000 25800 555024
rect 976 550000 1000 555000
rect 4000 550600 25800 555000
rect 27600 550600 61000 564000
rect 4000 550400 61000 550600
rect 65000 563700 320000 564000
rect 65000 563600 238200 563700
rect 65000 550400 126800 563600
rect 130800 558000 238200 563600
rect 239700 558000 320000 563700
rect 130800 557900 320000 558000
rect 130800 556400 263600 557900
rect 316600 556400 320000 557900
rect 130800 550400 320000 556400
rect 4000 550000 320000 550400
rect 976 549976 4024 550000
rect 198000 467800 200000 468000
rect 198000 466200 198200 467800
rect 199800 466200 200000 467800
rect 198000 466000 200000 466200
rect 122000 424200 152000 425400
rect 122000 419000 123600 424200
rect 30200 418600 123600 419000
rect 30200 409800 30600 418600
rect 39000 417800 123600 418600
rect 39000 416600 152000 417800
rect 39000 413600 123600 416600
rect 39000 412400 152000 413600
rect 39000 410600 123600 412400
rect 39000 409800 137600 410600
rect 30200 409400 137600 409800
rect 198000 361800 200000 362000
rect 198000 360200 198200 361800
rect 199800 360200 200000 361800
rect 198000 360000 200000 360200
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use BGR_lvs  BGR_lvs_0
timestamp 1669926749
transform 1 0 254230 0 1 568403
box -14230 -10403 62405 12600
use TX_line  TX_line_0
timestamp 1669931839
transform 1 0 200000 0 1 464000
box -24000 -130770 220000 24000
use VCO  VCO_0
timestamp 1663030914
transform 1 0 -7837 0 1 638742
box 31141 20430 65400 41673
use VCO  VCO_1
timestamp 1663030914
transform 0 1 115536 -1 0 464188
box 31141 20430 65400 41673
use VGA_routing  VGA_routing_0
timestamp 1667930445
transform 1 0 280 0 1 -18
box 165400 323622 584100 703354
<< labels >>
rlabel metal3 s 583520 269230 584800 269342 0 gpio_analog[0]
port 0 nsew signal bidirectional
rlabel metal3 s -800 381864 480 381976 0 gpio_analog[10]
port 1 nsew signal bidirectional
rlabel metal3 s -800 338642 480 338754 0 gpio_analog[11]
port 2 nsew signal bidirectional
rlabel metal3 s -800 295420 480 295532 0 gpio_analog[12]
port 3 nsew signal bidirectional
rlabel metal3 s -800 252398 480 252510 0 gpio_analog[13]
port 4 nsew signal bidirectional
rlabel metal3 s -800 124776 480 124888 0 gpio_analog[14]
port 5 nsew signal bidirectional
rlabel metal3 s -800 81554 480 81666 0 gpio_analog[15]
port 6 nsew signal bidirectional
rlabel metal3 s -800 38332 480 38444 0 gpio_analog[16]
port 7 nsew signal bidirectional
rlabel metal3 s -800 16910 480 17022 0 gpio_analog[17]
port 8 nsew signal bidirectional
rlabel metal3 s 583520 313652 584800 313764 0 gpio_analog[1]
port 9 nsew signal bidirectional
rlabel metal3 s 583520 358874 584800 358986 0 gpio_analog[2]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 405296 584800 405408 0 gpio_analog[3]
port 11 nsew signal bidirectional
rlabel metal3 s 583520 449718 584800 449830 0 gpio_analog[4]
port 12 nsew signal bidirectional
rlabel metal3 s 583520 494140 584800 494252 0 gpio_analog[5]
port 13 nsew signal bidirectional
rlabel metal3 s 583520 583562 584800 583674 0 gpio_analog[6]
port 14 nsew signal bidirectional
rlabel metal3 s -800 511530 480 511642 0 gpio_analog[7]
port 15 nsew signal bidirectional
rlabel metal3 s -800 468308 480 468420 0 gpio_analog[8]
port 16 nsew signal bidirectional
rlabel metal3 s -800 425086 480 425198 0 gpio_analog[9]
port 17 nsew signal bidirectional
rlabel metal3 s 583520 270412 584800 270524 0 gpio_noesd[0]
port 18 nsew signal bidirectional
rlabel metal3 s -800 380682 480 380794 0 gpio_noesd[10]
port 19 nsew signal bidirectional
rlabel metal3 s -800 337460 480 337572 0 gpio_noesd[11]
port 20 nsew signal bidirectional
rlabel metal3 s -800 294238 480 294350 0 gpio_noesd[12]
port 21 nsew signal bidirectional
rlabel metal3 s -800 251216 480 251328 0 gpio_noesd[13]
port 22 nsew signal bidirectional
rlabel metal3 s -800 123594 480 123706 0 gpio_noesd[14]
port 23 nsew signal bidirectional
rlabel metal3 s -800 80372 480 80484 0 gpio_noesd[15]
port 24 nsew signal bidirectional
rlabel metal3 s -800 37150 480 37262 0 gpio_noesd[16]
port 25 nsew signal bidirectional
rlabel metal3 s -800 15728 480 15840 0 gpio_noesd[17]
port 26 nsew signal bidirectional
rlabel metal3 s 583520 314834 584800 314946 0 gpio_noesd[1]
port 27 nsew signal bidirectional
rlabel metal3 s 583520 360056 584800 360168 0 gpio_noesd[2]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 406478 584800 406590 0 gpio_noesd[3]
port 29 nsew signal bidirectional
rlabel metal3 s 583520 450900 584800 451012 0 gpio_noesd[4]
port 30 nsew signal bidirectional
rlabel metal3 s 583520 495322 584800 495434 0 gpio_noesd[5]
port 31 nsew signal bidirectional
rlabel metal3 s 583520 584744 584800 584856 0 gpio_noesd[6]
port 32 nsew signal bidirectional
rlabel metal3 s -800 510348 480 510460 0 gpio_noesd[7]
port 33 nsew signal bidirectional
rlabel metal3 s -800 467126 480 467238 0 gpio_noesd[8]
port 34 nsew signal bidirectional
rlabel metal3 s -800 423904 480 424016 0 gpio_noesd[9]
port 35 nsew signal bidirectional
rlabel metal3 s 582300 677984 584800 682984 0 io_analog[0]
port 36 nsew signal bidirectional
rlabel metal3 0 680242 1700 685242 0 io_analog[10]
port 678 nsew
rlabel metal3 s 566594 702300 571594 704800 0 io_analog[1]
port 38 nsew signal bidirectional
rlabel metal3 s 465394 702300 470394 704800 0 io_analog[2]
port 39 nsew signal bidirectional
rlabel metal3 s 413394 702300 418394 704800 0 io_analog[3]
port 40 nsew signal bidirectional
rlabel metal3 s 329294 702300 334294 704800 0 io_analog[4]
port 41 nsew signal bidirectional
rlabel metal4 s 329294 702300 334294 704800 0 io_analog[4]
port 41 nsew signal bidirectional
rlabel metal5 s 329294 702300 334294 704800 0 io_analog[4]
port 41 nsew signal bidirectional
rlabel metal3 s 227594 702300 232594 704800 0 io_analog[5]
port 42 nsew signal bidirectional
rlabel metal4 s 227594 702300 232594 704800 0 io_analog[5]
port 42 nsew signal bidirectional
rlabel metal5 s 227594 702300 232594 704800 0 io_analog[5]
port 42 nsew signal bidirectional
rlabel metal3 s 175894 702300 180894 704800 0 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal4 s 175894 702300 180894 704800 0 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal5 s 175894 702300 180894 704800 0 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal3 s 120194 702300 125194 704800 0 io_analog[7]
port 44 nsew signal bidirectional
rlabel metal3 s 68194 702300 73194 704800 0 io_analog[8]
port 45 nsew signal bidirectional
rlabel metal3 s 16194 702300 21194 704800 0 io_analog[9]
port 46 nsew signal bidirectional
rlabel metal3 s 318994 702300 323994 704800 0 io_analog[4]
port 47 nsew signal bidirectional
rlabel metal4 s 318994 702300 323994 704800 0 io_analog[4]
port 47 nsew signal bidirectional
rlabel metal5 s 318994 702300 323994 704800 0 io_analog[4]
port 47 nsew signal bidirectional
rlabel metal3 s 217294 702300 222294 704800 0 io_analog[5]
port 48 nsew signal bidirectional
rlabel metal4 s 217294 702300 222294 704800 0 io_analog[5]
port 48 nsew signal bidirectional
rlabel metal5 s 217294 702300 222294 704800 0 io_analog[5]
port 48 nsew signal bidirectional
rlabel metal3 s 165594 702300 170594 704800 0 io_analog[6]
port 49 nsew signal bidirectional
rlabel metal4 s 165594 702300 170594 704800 0 io_analog[6]
port 49 nsew signal bidirectional
rlabel metal5 s 165594 702300 170594 704800 0 io_analog[6]
port 49 nsew signal bidirectional
rlabel metal3 s 326794 702300 328994 704800 0 io_clamp_high[0]
port 50 nsew signal bidirectional
rlabel metal3 s 225094 702300 227294 704800 0 io_clamp_high[1]
port 51 nsew signal bidirectional
rlabel metal3 s 173394 702300 175594 704800 0 io_clamp_high[2]
port 52 nsew signal bidirectional
rlabel metal3 s 324294 702300 326494 704800 0 io_clamp_low[0]
port 53 nsew signal bidirectional
rlabel metal3 s 222594 702300 224794 704800 0 io_clamp_low[1]
port 54 nsew signal bidirectional
rlabel metal3 s 170894 702300 173094 704800 0 io_clamp_low[2]
port 55 nsew signal bidirectional
rlabel metal3 s 583520 2726 584800 2838 0 io_in[0]
port 56 nsew signal input
rlabel metal3 s 583520 408842 584800 408954 0 io_in[10]
port 57 nsew signal input
rlabel metal3 s 583520 453264 584800 453376 0 io_in[11]
port 58 nsew signal input
rlabel metal3 s 583520 497686 584800 497798 0 io_in[12]
port 59 nsew signal input
rlabel metal3 s 583520 587108 584800 587220 0 io_in[13]
port 60 nsew signal input
rlabel metal3 s -800 507984 480 508096 0 io_in[14]
port 61 nsew signal input
rlabel metal3 s -800 464762 480 464874 0 io_in[15]
port 62 nsew signal input
rlabel metal3 s -800 421540 480 421652 0 io_in[16]
port 63 nsew signal input
rlabel metal3 s -800 378318 480 378430 0 io_in[17]
port 64 nsew signal input
rlabel metal3 s -800 335096 480 335208 0 io_in[18]
port 65 nsew signal input
rlabel metal3 s -800 291874 480 291986 0 io_in[19]
port 66 nsew signal input
rlabel metal3 s 583520 7454 584800 7566 0 io_in[1]
port 67 nsew signal input
rlabel metal3 s -800 248852 480 248964 0 io_in[20]
port 68 nsew signal input
rlabel metal3 s -800 121230 480 121342 0 io_in[21]
port 69 nsew signal input
rlabel metal3 s -800 78008 480 78120 0 io_in[22]
port 70 nsew signal input
rlabel metal3 s -800 34786 480 34898 0 io_in[23]
port 71 nsew signal input
rlabel metal3 s -800 13364 480 13476 0 io_in[24]
port 72 nsew signal input
rlabel metal3 s -800 8636 480 8748 0 io_in[25]
port 73 nsew signal input
rlabel metal3 s -800 3908 480 4020 0 io_in[26]
port 74 nsew signal input
rlabel metal3 s 583520 12182 584800 12294 0 io_in[2]
port 75 nsew signal input
rlabel metal3 s 583520 16910 584800 17022 0 io_in[3]
port 76 nsew signal input
rlabel metal3 s 583520 21638 584800 21750 0 io_in[4]
port 77 nsew signal input
rlabel metal3 s 583520 48096 584800 48208 0 io_in[5]
port 78 nsew signal input
rlabel metal3 s 583520 92754 584800 92866 0 io_in[6]
port 79 nsew signal input
rlabel metal3 s 583520 272776 584800 272888 0 io_in[7]
port 80 nsew signal input
rlabel metal3 s 583520 317198 584800 317310 0 io_in[8]
port 81 nsew signal input
rlabel metal3 s 583520 362420 584800 362532 0 io_in[9]
port 82 nsew signal input
rlabel metal3 s 583520 1544 584800 1656 0 io_in_3v3[0]
port 83 nsew signal input
rlabel metal3 s 583520 407660 584800 407772 0 io_in_3v3[10]
port 84 nsew signal input
rlabel metal3 s 583520 452082 584800 452194 0 io_in_3v3[11]
port 85 nsew signal input
rlabel metal3 s 583520 496504 584800 496616 0 io_in_3v3[12]
port 86 nsew signal input
rlabel metal3 s 583520 585926 584800 586038 0 io_in_3v3[13]
port 87 nsew signal input
rlabel metal3 s -800 509166 480 509278 0 io_in_3v3[14]
port 88 nsew signal input
rlabel metal3 s -800 465944 480 466056 0 io_in_3v3[15]
port 89 nsew signal input
rlabel metal3 s -800 422722 480 422834 0 io_in_3v3[16]
port 90 nsew signal input
rlabel metal3 s -800 379500 480 379612 0 io_in_3v3[17]
port 91 nsew signal input
rlabel metal3 s -800 336278 480 336390 0 io_in_3v3[18]
port 92 nsew signal input
rlabel metal3 s -800 293056 480 293168 0 io_in_3v3[19]
port 93 nsew signal input
rlabel metal3 s 583520 6272 584800 6384 0 io_in_3v3[1]
port 94 nsew signal input
rlabel metal3 s -800 250034 480 250146 0 io_in_3v3[20]
port 95 nsew signal input
rlabel metal3 s -800 122412 480 122524 0 io_in_3v3[21]
port 96 nsew signal input
rlabel metal3 s -800 79190 480 79302 0 io_in_3v3[22]
port 97 nsew signal input
rlabel metal3 s -800 35968 480 36080 0 io_in_3v3[23]
port 98 nsew signal input
rlabel metal3 s -800 14546 480 14658 0 io_in_3v3[24]
port 99 nsew signal input
rlabel metal3 s -800 9818 480 9930 0 io_in_3v3[25]
port 100 nsew signal input
rlabel metal3 s -800 5090 480 5202 0 io_in_3v3[26]
port 101 nsew signal input
rlabel metal3 s 583520 11000 584800 11112 0 io_in_3v3[2]
port 102 nsew signal input
rlabel metal3 s 583520 15728 584800 15840 0 io_in_3v3[3]
port 103 nsew signal input
rlabel metal3 s 583520 20456 584800 20568 0 io_in_3v3[4]
port 104 nsew signal input
rlabel metal3 s 583520 46914 584800 47026 0 io_in_3v3[5]
port 105 nsew signal input
rlabel metal3 s 583520 91572 584800 91684 0 io_in_3v3[6]
port 106 nsew signal input
rlabel metal3 s 583520 271594 584800 271706 0 io_in_3v3[7]
port 107 nsew signal input
rlabel metal3 s 583520 316016 584800 316128 0 io_in_3v3[8]
port 108 nsew signal input
rlabel metal3 s 583520 361238 584800 361350 0 io_in_3v3[9]
port 109 nsew signal input
rlabel metal3 s 583520 5090 584800 5202 0 io_oeb[0]
port 110 nsew signal tristate
rlabel metal3 s 583520 411206 584800 411318 0 io_oeb[10]
port 111 nsew signal tristate
rlabel metal3 s 583520 455628 584800 455740 0 io_oeb[11]
port 112 nsew signal tristate
rlabel metal3 s 583520 500050 584800 500162 0 io_oeb[12]
port 113 nsew signal tristate
rlabel metal3 s 583520 589472 584800 589584 0 io_oeb[13]
port 114 nsew signal tristate
rlabel metal3 s -800 505620 480 505732 0 io_oeb[14]
port 115 nsew signal tristate
rlabel metal3 s -800 462398 480 462510 0 io_oeb[15]
port 116 nsew signal tristate
rlabel metal3 s -800 419176 480 419288 0 io_oeb[16]
port 117 nsew signal tristate
rlabel metal3 s -800 375954 480 376066 0 io_oeb[17]
port 118 nsew signal tristate
rlabel metal3 s -800 332732 480 332844 0 io_oeb[18]
port 119 nsew signal tristate
rlabel metal3 s -800 289510 480 289622 0 io_oeb[19]
port 120 nsew signal tristate
rlabel metal3 s 583520 9818 584800 9930 0 io_oeb[1]
port 121 nsew signal tristate
rlabel metal3 s -800 246488 480 246600 0 io_oeb[20]
port 122 nsew signal tristate
rlabel metal3 s -800 118866 480 118978 0 io_oeb[21]
port 123 nsew signal tristate
rlabel metal3 s -800 75644 480 75756 0 io_oeb[22]
port 124 nsew signal tristate
rlabel metal3 s -800 32422 480 32534 0 io_oeb[23]
port 125 nsew signal tristate
rlabel metal3 s -800 11000 480 11112 0 io_oeb[24]
port 126 nsew signal tristate
rlabel metal3 s -800 6272 480 6384 0 io_oeb[25]
port 127 nsew signal tristate
rlabel metal3 s -800 1544 480 1656 0 io_oeb[26]
port 128 nsew signal tristate
rlabel metal3 s 583520 14546 584800 14658 0 io_oeb[2]
port 129 nsew signal tristate
rlabel metal3 s 583520 19274 584800 19386 0 io_oeb[3]
port 130 nsew signal tristate
rlabel metal3 s 583520 24002 584800 24114 0 io_oeb[4]
port 131 nsew signal tristate
rlabel metal3 s 583520 50460 584800 50572 0 io_oeb[5]
port 132 nsew signal tristate
rlabel metal3 s 583520 95118 584800 95230 0 io_oeb[6]
port 133 nsew signal tristate
rlabel metal3 s 583520 275140 584800 275252 0 io_oeb[7]
port 134 nsew signal tristate
rlabel metal3 s 583520 319562 584800 319674 0 io_oeb[8]
port 135 nsew signal tristate
rlabel metal3 s 583520 364784 584800 364896 0 io_oeb[9]
port 136 nsew signal tristate
rlabel metal3 s 583520 3908 584800 4020 0 io_out[0]
port 137 nsew signal tristate
rlabel metal3 s 583520 410024 584800 410136 0 io_out[10]
port 138 nsew signal tristate
rlabel metal3 s 583520 454446 584800 454558 0 io_out[11]
port 139 nsew signal tristate
rlabel metal3 s 583520 498868 584800 498980 0 io_out[12]
port 140 nsew signal tristate
rlabel metal3 s 583520 588290 584800 588402 0 io_out[13]
port 141 nsew signal tristate
rlabel metal3 s -800 506802 480 506914 0 io_out[14]
port 142 nsew signal tristate
rlabel metal3 s -800 463580 480 463692 0 io_out[15]
port 143 nsew signal tristate
rlabel metal3 s -800 420358 480 420470 0 io_out[16]
port 144 nsew signal tristate
rlabel metal3 s -800 377136 480 377248 0 io_out[17]
port 145 nsew signal tristate
rlabel metal3 s -800 333914 480 334026 0 io_out[18]
port 146 nsew signal tristate
rlabel metal3 s -800 290692 480 290804 0 io_out[19]
port 147 nsew signal tristate
rlabel metal3 s 583520 8636 584800 8748 0 io_out[1]
port 148 nsew signal tristate
rlabel metal3 s -800 247670 480 247782 0 io_out[20]
port 149 nsew signal tristate
rlabel metal3 s -800 120048 480 120160 0 io_out[21]
port 150 nsew signal tristate
rlabel metal3 s -800 76826 480 76938 0 io_out[22]
port 151 nsew signal tristate
rlabel metal3 s -800 33604 480 33716 0 io_out[23]
port 152 nsew signal tristate
rlabel metal3 s -800 12182 480 12294 0 io_out[24]
port 153 nsew signal tristate
rlabel metal3 s -800 7454 480 7566 0 io_out[25]
port 154 nsew signal tristate
rlabel metal3 s -800 2726 480 2838 0 io_out[26]
port 155 nsew signal tristate
rlabel metal3 s 583520 13364 584800 13476 0 io_out[2]
port 156 nsew signal tristate
rlabel metal3 s 583520 18092 584800 18204 0 io_out[3]
port 157 nsew signal tristate
rlabel metal3 s 583520 22820 584800 22932 0 io_out[4]
port 158 nsew signal tristate
rlabel metal3 s 583520 49278 584800 49390 0 io_out[5]
port 159 nsew signal tristate
rlabel metal3 s 583520 93936 584800 94048 0 io_out[6]
port 160 nsew signal tristate
rlabel metal3 s 583520 273958 584800 274070 0 io_out[7]
port 161 nsew signal tristate
rlabel metal3 s 583520 318380 584800 318492 0 io_out[8]
port 162 nsew signal tristate
rlabel metal3 s 583520 363602 584800 363714 0 io_out[9]
port 163 nsew signal tristate
rlabel metal2 s 125816 -800 125928 480 0 la_data_in[0]
port 164 nsew signal input
rlabel metal2 s 480416 -800 480528 480 0 la_data_in[100]
port 165 nsew signal input
rlabel metal2 s 483962 -800 484074 480 0 la_data_in[101]
port 166 nsew signal input
rlabel metal2 s 487508 -800 487620 480 0 la_data_in[102]
port 167 nsew signal input
rlabel metal2 s 491054 -800 491166 480 0 la_data_in[103]
port 168 nsew signal input
rlabel metal2 s 494600 -800 494712 480 0 la_data_in[104]
port 169 nsew signal input
rlabel metal2 s 498146 -800 498258 480 0 la_data_in[105]
port 170 nsew signal input
rlabel metal2 s 501692 -800 501804 480 0 la_data_in[106]
port 171 nsew signal input
rlabel metal2 s 505238 -800 505350 480 0 la_data_in[107]
port 172 nsew signal input
rlabel metal2 s 508784 -800 508896 480 0 la_data_in[108]
port 173 nsew signal input
rlabel metal2 s 512330 -800 512442 480 0 la_data_in[109]
port 174 nsew signal input
rlabel metal2 s 161276 -800 161388 480 0 la_data_in[10]
port 175 nsew signal input
rlabel metal2 s 515876 -800 515988 480 0 la_data_in[110]
port 176 nsew signal input
rlabel metal2 s 519422 -800 519534 480 0 la_data_in[111]
port 177 nsew signal input
rlabel metal2 s 522968 -800 523080 480 0 la_data_in[112]
port 178 nsew signal input
rlabel metal2 s 526514 -800 526626 480 0 la_data_in[113]
port 179 nsew signal input
rlabel metal2 s 530060 -800 530172 480 0 la_data_in[114]
port 180 nsew signal input
rlabel metal2 s 533606 -800 533718 480 0 la_data_in[115]
port 181 nsew signal input
rlabel metal2 s 537152 -800 537264 480 0 la_data_in[116]
port 182 nsew signal input
rlabel metal2 s 540698 -800 540810 480 0 la_data_in[117]
port 183 nsew signal input
rlabel metal2 s 544244 -800 544356 480 0 la_data_in[118]
port 184 nsew signal input
rlabel metal2 s 547790 -800 547902 480 0 la_data_in[119]
port 185 nsew signal input
rlabel metal2 s 164822 -800 164934 480 0 la_data_in[11]
port 186 nsew signal input
rlabel metal2 s 551336 -800 551448 480 0 la_data_in[120]
port 187 nsew signal input
rlabel metal2 s 554882 -800 554994 480 0 la_data_in[121]
port 188 nsew signal input
rlabel metal2 s 558428 -800 558540 480 0 la_data_in[122]
port 189 nsew signal input
rlabel metal2 s 561974 -800 562086 480 0 la_data_in[123]
port 190 nsew signal input
rlabel metal2 s 565520 -800 565632 480 0 la_data_in[124]
port 191 nsew signal input
rlabel metal2 s 569066 -800 569178 480 0 la_data_in[125]
port 192 nsew signal input
rlabel metal2 s 572612 -800 572724 480 0 la_data_in[126]
port 193 nsew signal input
rlabel metal2 s 576158 -800 576270 480 0 la_data_in[127]
port 194 nsew signal input
rlabel metal2 s 168368 -800 168480 480 0 la_data_in[12]
port 195 nsew signal input
rlabel metal2 s 171914 -800 172026 480 0 la_data_in[13]
port 196 nsew signal input
rlabel metal2 s 175460 -800 175572 480 0 la_data_in[14]
port 197 nsew signal input
rlabel metal2 s 179006 -800 179118 480 0 la_data_in[15]
port 198 nsew signal input
rlabel metal2 s 182552 -800 182664 480 0 la_data_in[16]
port 199 nsew signal input
rlabel metal2 s 186098 -800 186210 480 0 la_data_in[17]
port 200 nsew signal input
rlabel metal2 s 189644 -800 189756 480 0 la_data_in[18]
port 201 nsew signal input
rlabel metal2 s 193190 -800 193302 480 0 la_data_in[19]
port 202 nsew signal input
rlabel metal2 s 129362 -800 129474 480 0 la_data_in[1]
port 203 nsew signal input
rlabel metal2 s 196736 -800 196848 480 0 la_data_in[20]
port 204 nsew signal input
rlabel metal2 s 200282 -800 200394 480 0 la_data_in[21]
port 205 nsew signal input
rlabel metal2 s 203828 -800 203940 480 0 la_data_in[22]
port 206 nsew signal input
rlabel metal2 s 207374 -800 207486 480 0 la_data_in[23]
port 207 nsew signal input
rlabel metal2 s 210920 -800 211032 480 0 la_data_in[24]
port 208 nsew signal input
rlabel metal2 s 214466 -800 214578 480 0 la_data_in[25]
port 209 nsew signal input
rlabel metal2 s 218012 -800 218124 480 0 la_data_in[26]
port 210 nsew signal input
rlabel metal2 s 221558 -800 221670 480 0 la_data_in[27]
port 211 nsew signal input
rlabel metal2 s 225104 -800 225216 480 0 la_data_in[28]
port 212 nsew signal input
rlabel metal2 s 228650 -800 228762 480 0 la_data_in[29]
port 213 nsew signal input
rlabel metal2 s 132908 -800 133020 480 0 la_data_in[2]
port 214 nsew signal input
rlabel metal2 s 232196 -800 232308 480 0 la_data_in[30]
port 215 nsew signal input
rlabel metal2 s 235742 -800 235854 480 0 la_data_in[31]
port 216 nsew signal input
rlabel metal2 s 239288 -800 239400 480 0 la_data_in[32]
port 217 nsew signal input
rlabel metal2 s 242834 -800 242946 480 0 la_data_in[33]
port 218 nsew signal input
rlabel metal2 s 246380 -800 246492 480 0 la_data_in[34]
port 219 nsew signal input
rlabel metal2 s 249926 -800 250038 480 0 la_data_in[35]
port 220 nsew signal input
rlabel metal2 s 253472 -800 253584 480 0 la_data_in[36]
port 221 nsew signal input
rlabel metal2 s 257018 -800 257130 480 0 la_data_in[37]
port 222 nsew signal input
rlabel metal2 s 260564 -800 260676 480 0 la_data_in[38]
port 223 nsew signal input
rlabel metal2 s 264110 -800 264222 480 0 la_data_in[39]
port 224 nsew signal input
rlabel metal2 s 136454 -800 136566 480 0 la_data_in[3]
port 225 nsew signal input
rlabel metal2 s 267656 -800 267768 480 0 la_data_in[40]
port 226 nsew signal input
rlabel metal2 s 271202 -800 271314 480 0 la_data_in[41]
port 227 nsew signal input
rlabel metal2 s 274748 -800 274860 480 0 la_data_in[42]
port 228 nsew signal input
rlabel metal2 s 278294 -800 278406 480 0 la_data_in[43]
port 229 nsew signal input
rlabel metal2 s 281840 -800 281952 480 0 la_data_in[44]
port 230 nsew signal input
rlabel metal2 s 285386 -800 285498 480 0 la_data_in[45]
port 231 nsew signal input
rlabel metal2 s 288932 -800 289044 480 0 la_data_in[46]
port 232 nsew signal input
rlabel metal2 s 292478 -800 292590 480 0 la_data_in[47]
port 233 nsew signal input
rlabel metal2 s 296024 -800 296136 480 0 la_data_in[48]
port 234 nsew signal input
rlabel metal2 s 299570 -800 299682 480 0 la_data_in[49]
port 235 nsew signal input
rlabel metal2 s 140000 -800 140112 480 0 la_data_in[4]
port 236 nsew signal input
rlabel metal2 s 303116 -800 303228 480 0 la_data_in[50]
port 237 nsew signal input
rlabel metal2 s 306662 -800 306774 480 0 la_data_in[51]
port 238 nsew signal input
rlabel metal2 s 310208 -800 310320 480 0 la_data_in[52]
port 239 nsew signal input
rlabel metal2 s 313754 -800 313866 480 0 la_data_in[53]
port 240 nsew signal input
rlabel metal2 s 317300 -800 317412 480 0 la_data_in[54]
port 241 nsew signal input
rlabel metal2 s 320846 -800 320958 480 0 la_data_in[55]
port 242 nsew signal input
rlabel metal2 s 324392 -800 324504 480 0 la_data_in[56]
port 243 nsew signal input
rlabel metal2 s 327938 -800 328050 480 0 la_data_in[57]
port 244 nsew signal input
rlabel metal2 s 331484 -800 331596 480 0 la_data_in[58]
port 245 nsew signal input
rlabel metal2 s 335030 -800 335142 480 0 la_data_in[59]
port 246 nsew signal input
rlabel metal2 s 143546 -800 143658 480 0 la_data_in[5]
port 247 nsew signal input
rlabel metal2 s 338576 -800 338688 480 0 la_data_in[60]
port 248 nsew signal input
rlabel metal2 s 342122 -800 342234 480 0 la_data_in[61]
port 249 nsew signal input
rlabel metal2 s 345668 -800 345780 480 0 la_data_in[62]
port 250 nsew signal input
rlabel metal2 s 349214 -800 349326 480 0 la_data_in[63]
port 251 nsew signal input
rlabel metal2 s 352760 -800 352872 480 0 la_data_in[64]
port 252 nsew signal input
rlabel metal2 s 356306 -800 356418 480 0 la_data_in[65]
port 253 nsew signal input
rlabel metal2 s 359852 -800 359964 480 0 la_data_in[66]
port 254 nsew signal input
rlabel metal2 s 363398 -800 363510 480 0 la_data_in[67]
port 255 nsew signal input
rlabel metal2 s 366944 -800 367056 480 0 la_data_in[68]
port 256 nsew signal input
rlabel metal2 s 370490 -800 370602 480 0 la_data_in[69]
port 257 nsew signal input
rlabel metal2 s 147092 -800 147204 480 0 la_data_in[6]
port 258 nsew signal input
rlabel metal2 s 374036 -800 374148 480 0 la_data_in[70]
port 259 nsew signal input
rlabel metal2 s 377582 -800 377694 480 0 la_data_in[71]
port 260 nsew signal input
rlabel metal2 s 381128 -800 381240 480 0 la_data_in[72]
port 261 nsew signal input
rlabel metal2 s 384674 -800 384786 480 0 la_data_in[73]
port 262 nsew signal input
rlabel metal2 s 388220 -800 388332 480 0 la_data_in[74]
port 263 nsew signal input
rlabel metal2 s 391766 -800 391878 480 0 la_data_in[75]
port 264 nsew signal input
rlabel metal2 s 395312 -800 395424 480 0 la_data_in[76]
port 265 nsew signal input
rlabel metal2 s 398858 -800 398970 480 0 la_data_in[77]
port 266 nsew signal input
rlabel metal2 s 402404 -800 402516 480 0 la_data_in[78]
port 267 nsew signal input
rlabel metal2 s 405950 -800 406062 480 0 la_data_in[79]
port 268 nsew signal input
rlabel metal2 s 150638 -800 150750 480 0 la_data_in[7]
port 269 nsew signal input
rlabel metal2 s 409496 -800 409608 480 0 la_data_in[80]
port 270 nsew signal input
rlabel metal2 s 413042 -800 413154 480 0 la_data_in[81]
port 271 nsew signal input
rlabel metal2 s 416588 -800 416700 480 0 la_data_in[82]
port 272 nsew signal input
rlabel metal2 s 420134 -800 420246 480 0 la_data_in[83]
port 273 nsew signal input
rlabel metal2 s 423680 -800 423792 480 0 la_data_in[84]
port 274 nsew signal input
rlabel metal2 s 427226 -800 427338 480 0 la_data_in[85]
port 275 nsew signal input
rlabel metal2 s 430772 -800 430884 480 0 la_data_in[86]
port 276 nsew signal input
rlabel metal2 s 434318 -800 434430 480 0 la_data_in[87]
port 277 nsew signal input
rlabel metal2 s 437864 -800 437976 480 0 la_data_in[88]
port 278 nsew signal input
rlabel metal2 s 441410 -800 441522 480 0 la_data_in[89]
port 279 nsew signal input
rlabel metal2 s 154184 -800 154296 480 0 la_data_in[8]
port 280 nsew signal input
rlabel metal2 s 444956 -800 445068 480 0 la_data_in[90]
port 281 nsew signal input
rlabel metal2 s 448502 -800 448614 480 0 la_data_in[91]
port 282 nsew signal input
rlabel metal2 s 452048 -800 452160 480 0 la_data_in[92]
port 283 nsew signal input
rlabel metal2 s 455594 -800 455706 480 0 la_data_in[93]
port 284 nsew signal input
rlabel metal2 s 459140 -800 459252 480 0 la_data_in[94]
port 285 nsew signal input
rlabel metal2 s 462686 -800 462798 480 0 la_data_in[95]
port 286 nsew signal input
rlabel metal2 s 466232 -800 466344 480 0 la_data_in[96]
port 287 nsew signal input
rlabel metal2 s 469778 -800 469890 480 0 la_data_in[97]
port 288 nsew signal input
rlabel metal2 s 473324 -800 473436 480 0 la_data_in[98]
port 289 nsew signal input
rlabel metal2 s 476870 -800 476982 480 0 la_data_in[99]
port 290 nsew signal input
rlabel metal2 s 157730 -800 157842 480 0 la_data_in[9]
port 291 nsew signal input
rlabel metal2 s 126998 -800 127110 480 0 la_data_out[0]
port 292 nsew signal tristate
rlabel metal2 s 481598 -800 481710 480 0 la_data_out[100]
port 293 nsew signal tristate
rlabel metal2 s 485144 -800 485256 480 0 la_data_out[101]
port 294 nsew signal tristate
rlabel metal2 s 488690 -800 488802 480 0 la_data_out[102]
port 295 nsew signal tristate
rlabel metal2 s 492236 -800 492348 480 0 la_data_out[103]
port 296 nsew signal tristate
rlabel metal2 s 495782 -800 495894 480 0 la_data_out[104]
port 297 nsew signal tristate
rlabel metal2 s 499328 -800 499440 480 0 la_data_out[105]
port 298 nsew signal tristate
rlabel metal2 s 502874 -800 502986 480 0 la_data_out[106]
port 299 nsew signal tristate
rlabel metal2 s 506420 -800 506532 480 0 la_data_out[107]
port 300 nsew signal tristate
rlabel metal2 s 509966 -800 510078 480 0 la_data_out[108]
port 301 nsew signal tristate
rlabel metal2 s 513512 -800 513624 480 0 la_data_out[109]
port 302 nsew signal tristate
rlabel metal2 s 162458 -800 162570 480 0 la_data_out[10]
port 303 nsew signal tristate
rlabel metal2 s 517058 -800 517170 480 0 la_data_out[110]
port 304 nsew signal tristate
rlabel metal2 s 520604 -800 520716 480 0 la_data_out[111]
port 305 nsew signal tristate
rlabel metal2 s 524150 -800 524262 480 0 la_data_out[112]
port 306 nsew signal tristate
rlabel metal2 s 527696 -800 527808 480 0 la_data_out[113]
port 307 nsew signal tristate
rlabel metal2 s 531242 -800 531354 480 0 la_data_out[114]
port 308 nsew signal tristate
rlabel metal2 s 534788 -800 534900 480 0 la_data_out[115]
port 309 nsew signal tristate
rlabel metal2 s 538334 -800 538446 480 0 la_data_out[116]
port 310 nsew signal tristate
rlabel metal2 s 541880 -800 541992 480 0 la_data_out[117]
port 311 nsew signal tristate
rlabel metal2 s 545426 -800 545538 480 0 la_data_out[118]
port 312 nsew signal tristate
rlabel metal2 s 548972 -800 549084 480 0 la_data_out[119]
port 313 nsew signal tristate
rlabel metal2 s 166004 -800 166116 480 0 la_data_out[11]
port 314 nsew signal tristate
rlabel metal2 s 552518 -800 552630 480 0 la_data_out[120]
port 315 nsew signal tristate
rlabel metal2 s 556064 -800 556176 480 0 la_data_out[121]
port 316 nsew signal tristate
rlabel metal2 s 559610 -800 559722 480 0 la_data_out[122]
port 317 nsew signal tristate
rlabel metal2 s 563156 -800 563268 480 0 la_data_out[123]
port 318 nsew signal tristate
rlabel metal2 s 566702 -800 566814 480 0 la_data_out[124]
port 319 nsew signal tristate
rlabel metal2 s 570248 -800 570360 480 0 la_data_out[125]
port 320 nsew signal tristate
rlabel metal2 s 573794 -800 573906 480 0 la_data_out[126]
port 321 nsew signal tristate
rlabel metal2 s 577340 -800 577452 480 0 la_data_out[127]
port 322 nsew signal tristate
rlabel metal2 s 169550 -800 169662 480 0 la_data_out[12]
port 323 nsew signal tristate
rlabel metal2 s 173096 -800 173208 480 0 la_data_out[13]
port 324 nsew signal tristate
rlabel metal2 s 176642 -800 176754 480 0 la_data_out[14]
port 325 nsew signal tristate
rlabel metal2 s 180188 -800 180300 480 0 la_data_out[15]
port 326 nsew signal tristate
rlabel metal2 s 183734 -800 183846 480 0 la_data_out[16]
port 327 nsew signal tristate
rlabel metal2 s 187280 -800 187392 480 0 la_data_out[17]
port 328 nsew signal tristate
rlabel metal2 s 190826 -800 190938 480 0 la_data_out[18]
port 329 nsew signal tristate
rlabel metal2 s 194372 -800 194484 480 0 la_data_out[19]
port 330 nsew signal tristate
rlabel metal2 s 130544 -800 130656 480 0 la_data_out[1]
port 331 nsew signal tristate
rlabel metal2 s 197918 -800 198030 480 0 la_data_out[20]
port 332 nsew signal tristate
rlabel metal2 s 201464 -800 201576 480 0 la_data_out[21]
port 333 nsew signal tristate
rlabel metal2 s 205010 -800 205122 480 0 la_data_out[22]
port 334 nsew signal tristate
rlabel metal2 s 208556 -800 208668 480 0 la_data_out[23]
port 335 nsew signal tristate
rlabel metal2 s 212102 -800 212214 480 0 la_data_out[24]
port 336 nsew signal tristate
rlabel metal2 s 215648 -800 215760 480 0 la_data_out[25]
port 337 nsew signal tristate
rlabel metal2 s 219194 -800 219306 480 0 la_data_out[26]
port 338 nsew signal tristate
rlabel metal2 s 222740 -800 222852 480 0 la_data_out[27]
port 339 nsew signal tristate
rlabel metal2 s 226286 -800 226398 480 0 la_data_out[28]
port 340 nsew signal tristate
rlabel metal2 s 229832 -800 229944 480 0 la_data_out[29]
port 341 nsew signal tristate
rlabel metal2 s 134090 -800 134202 480 0 la_data_out[2]
port 342 nsew signal tristate
rlabel metal2 s 233378 -800 233490 480 0 la_data_out[30]
port 343 nsew signal tristate
rlabel metal2 s 236924 -800 237036 480 0 la_data_out[31]
port 344 nsew signal tristate
rlabel metal2 s 240470 -800 240582 480 0 la_data_out[32]
port 345 nsew signal tristate
rlabel metal2 s 244016 -800 244128 480 0 la_data_out[33]
port 346 nsew signal tristate
rlabel metal2 s 247562 -800 247674 480 0 la_data_out[34]
port 347 nsew signal tristate
rlabel metal2 s 251108 -800 251220 480 0 la_data_out[35]
port 348 nsew signal tristate
rlabel metal2 s 254654 -800 254766 480 0 la_data_out[36]
port 349 nsew signal tristate
rlabel metal2 s 258200 -800 258312 480 0 la_data_out[37]
port 350 nsew signal tristate
rlabel metal2 s 261746 -800 261858 480 0 la_data_out[38]
port 351 nsew signal tristate
rlabel metal2 s 265292 -800 265404 480 0 la_data_out[39]
port 352 nsew signal tristate
rlabel metal2 s 137636 -800 137748 480 0 la_data_out[3]
port 353 nsew signal tristate
rlabel metal2 s 268838 -800 268950 480 0 la_data_out[40]
port 354 nsew signal tristate
rlabel metal2 s 272384 -800 272496 480 0 la_data_out[41]
port 355 nsew signal tristate
rlabel metal2 s 275930 -800 276042 480 0 la_data_out[42]
port 356 nsew signal tristate
rlabel metal2 s 279476 -800 279588 480 0 la_data_out[43]
port 357 nsew signal tristate
rlabel metal2 s 283022 -800 283134 480 0 la_data_out[44]
port 358 nsew signal tristate
rlabel metal2 s 286568 -800 286680 480 0 la_data_out[45]
port 359 nsew signal tristate
rlabel metal2 s 290114 -800 290226 480 0 la_data_out[46]
port 360 nsew signal tristate
rlabel metal2 s 293660 -800 293772 480 0 la_data_out[47]
port 361 nsew signal tristate
rlabel metal2 s 297206 -800 297318 480 0 la_data_out[48]
port 362 nsew signal tristate
rlabel metal2 s 300752 -800 300864 480 0 la_data_out[49]
port 363 nsew signal tristate
rlabel metal2 s 141182 -800 141294 480 0 la_data_out[4]
port 364 nsew signal tristate
rlabel metal2 s 304298 -800 304410 480 0 la_data_out[50]
port 365 nsew signal tristate
rlabel metal2 s 307844 -800 307956 480 0 la_data_out[51]
port 366 nsew signal tristate
rlabel metal2 s 311390 -800 311502 480 0 la_data_out[52]
port 367 nsew signal tristate
rlabel metal2 s 314936 -800 315048 480 0 la_data_out[53]
port 368 nsew signal tristate
rlabel metal2 s 318482 -800 318594 480 0 la_data_out[54]
port 369 nsew signal tristate
rlabel metal2 s 322028 -800 322140 480 0 la_data_out[55]
port 370 nsew signal tristate
rlabel metal2 s 325574 -800 325686 480 0 la_data_out[56]
port 371 nsew signal tristate
rlabel metal2 s 329120 -800 329232 480 0 la_data_out[57]
port 372 nsew signal tristate
rlabel metal2 s 332666 -800 332778 480 0 la_data_out[58]
port 373 nsew signal tristate
rlabel metal2 s 336212 -800 336324 480 0 la_data_out[59]
port 374 nsew signal tristate
rlabel metal2 s 144728 -800 144840 480 0 la_data_out[5]
port 375 nsew signal tristate
rlabel metal2 s 339758 -800 339870 480 0 la_data_out[60]
port 376 nsew signal tristate
rlabel metal2 s 343304 -800 343416 480 0 la_data_out[61]
port 377 nsew signal tristate
rlabel metal2 s 346850 -800 346962 480 0 la_data_out[62]
port 378 nsew signal tristate
rlabel metal2 s 350396 -800 350508 480 0 la_data_out[63]
port 379 nsew signal tristate
rlabel metal2 s 353942 -800 354054 480 0 la_data_out[64]
port 380 nsew signal tristate
rlabel metal2 s 357488 -800 357600 480 0 la_data_out[65]
port 381 nsew signal tristate
rlabel metal2 s 361034 -800 361146 480 0 la_data_out[66]
port 382 nsew signal tristate
rlabel metal2 s 364580 -800 364692 480 0 la_data_out[67]
port 383 nsew signal tristate
rlabel metal2 s 368126 -800 368238 480 0 la_data_out[68]
port 384 nsew signal tristate
rlabel metal2 s 371672 -800 371784 480 0 la_data_out[69]
port 385 nsew signal tristate
rlabel metal2 s 148274 -800 148386 480 0 la_data_out[6]
port 386 nsew signal tristate
rlabel metal2 s 375218 -800 375330 480 0 la_data_out[70]
port 387 nsew signal tristate
rlabel metal2 s 378764 -800 378876 480 0 la_data_out[71]
port 388 nsew signal tristate
rlabel metal2 s 382310 -800 382422 480 0 la_data_out[72]
port 389 nsew signal tristate
rlabel metal2 s 385856 -800 385968 480 0 la_data_out[73]
port 390 nsew signal tristate
rlabel metal2 s 389402 -800 389514 480 0 la_data_out[74]
port 391 nsew signal tristate
rlabel metal2 s 392948 -800 393060 480 0 la_data_out[75]
port 392 nsew signal tristate
rlabel metal2 s 396494 -800 396606 480 0 la_data_out[76]
port 393 nsew signal tristate
rlabel metal2 s 400040 -800 400152 480 0 la_data_out[77]
port 394 nsew signal tristate
rlabel metal2 s 403586 -800 403698 480 0 la_data_out[78]
port 395 nsew signal tristate
rlabel metal2 s 407132 -800 407244 480 0 la_data_out[79]
port 396 nsew signal tristate
rlabel metal2 s 151820 -800 151932 480 0 la_data_out[7]
port 397 nsew signal tristate
rlabel metal2 s 410678 -800 410790 480 0 la_data_out[80]
port 398 nsew signal tristate
rlabel metal2 s 414224 -800 414336 480 0 la_data_out[81]
port 399 nsew signal tristate
rlabel metal2 s 417770 -800 417882 480 0 la_data_out[82]
port 400 nsew signal tristate
rlabel metal2 s 421316 -800 421428 480 0 la_data_out[83]
port 401 nsew signal tristate
rlabel metal2 s 424862 -800 424974 480 0 la_data_out[84]
port 402 nsew signal tristate
rlabel metal2 s 428408 -800 428520 480 0 la_data_out[85]
port 403 nsew signal tristate
rlabel metal2 s 431954 -800 432066 480 0 la_data_out[86]
port 404 nsew signal tristate
rlabel metal2 s 435500 -800 435612 480 0 la_data_out[87]
port 405 nsew signal tristate
rlabel metal2 s 439046 -800 439158 480 0 la_data_out[88]
port 406 nsew signal tristate
rlabel metal2 s 442592 -800 442704 480 0 la_data_out[89]
port 407 nsew signal tristate
rlabel metal2 s 155366 -800 155478 480 0 la_data_out[8]
port 408 nsew signal tristate
rlabel metal2 s 446138 -800 446250 480 0 la_data_out[90]
port 409 nsew signal tristate
rlabel metal2 s 449684 -800 449796 480 0 la_data_out[91]
port 410 nsew signal tristate
rlabel metal2 s 453230 -800 453342 480 0 la_data_out[92]
port 411 nsew signal tristate
rlabel metal2 s 456776 -800 456888 480 0 la_data_out[93]
port 412 nsew signal tristate
rlabel metal2 s 460322 -800 460434 480 0 la_data_out[94]
port 413 nsew signal tristate
rlabel metal2 s 463868 -800 463980 480 0 la_data_out[95]
port 414 nsew signal tristate
rlabel metal2 s 467414 -800 467526 480 0 la_data_out[96]
port 415 nsew signal tristate
rlabel metal2 s 470960 -800 471072 480 0 la_data_out[97]
port 416 nsew signal tristate
rlabel metal2 s 474506 -800 474618 480 0 la_data_out[98]
port 417 nsew signal tristate
rlabel metal2 s 478052 -800 478164 480 0 la_data_out[99]
port 418 nsew signal tristate
rlabel metal2 s 158912 -800 159024 480 0 la_data_out[9]
port 419 nsew signal tristate
rlabel metal2 s 128180 -800 128292 480 0 la_oenb[0]
port 420 nsew signal input
rlabel metal2 s 482780 -800 482892 480 0 la_oenb[100]
port 421 nsew signal input
rlabel metal2 s 486326 -800 486438 480 0 la_oenb[101]
port 422 nsew signal input
rlabel metal2 s 489872 -800 489984 480 0 la_oenb[102]
port 423 nsew signal input
rlabel metal2 s 493418 -800 493530 480 0 la_oenb[103]
port 424 nsew signal input
rlabel metal2 s 496964 -800 497076 480 0 la_oenb[104]
port 425 nsew signal input
rlabel metal2 s 500510 -800 500622 480 0 la_oenb[105]
port 426 nsew signal input
rlabel metal2 s 504056 -800 504168 480 0 la_oenb[106]
port 427 nsew signal input
rlabel metal2 s 507602 -800 507714 480 0 la_oenb[107]
port 428 nsew signal input
rlabel metal2 s 511148 -800 511260 480 0 la_oenb[108]
port 429 nsew signal input
rlabel metal2 s 514694 -800 514806 480 0 la_oenb[109]
port 430 nsew signal input
rlabel metal2 s 163640 -800 163752 480 0 la_oenb[10]
port 431 nsew signal input
rlabel metal2 s 518240 -800 518352 480 0 la_oenb[110]
port 432 nsew signal input
rlabel metal2 s 521786 -800 521898 480 0 la_oenb[111]
port 433 nsew signal input
rlabel metal2 s 525332 -800 525444 480 0 la_oenb[112]
port 434 nsew signal input
rlabel metal2 s 528878 -800 528990 480 0 la_oenb[113]
port 435 nsew signal input
rlabel metal2 s 532424 -800 532536 480 0 la_oenb[114]
port 436 nsew signal input
rlabel metal2 s 535970 -800 536082 480 0 la_oenb[115]
port 437 nsew signal input
rlabel metal2 s 539516 -800 539628 480 0 la_oenb[116]
port 438 nsew signal input
rlabel metal2 s 543062 -800 543174 480 0 la_oenb[117]
port 439 nsew signal input
rlabel metal2 s 546608 -800 546720 480 0 la_oenb[118]
port 440 nsew signal input
rlabel metal2 s 550154 -800 550266 480 0 la_oenb[119]
port 441 nsew signal input
rlabel metal2 s 167186 -800 167298 480 0 la_oenb[11]
port 442 nsew signal input
rlabel metal2 s 553700 -800 553812 480 0 la_oenb[120]
port 443 nsew signal input
rlabel metal2 s 557246 -800 557358 480 0 la_oenb[121]
port 444 nsew signal input
rlabel metal2 s 560792 -800 560904 480 0 la_oenb[122]
port 445 nsew signal input
rlabel metal2 s 564338 -800 564450 480 0 la_oenb[123]
port 446 nsew signal input
rlabel metal2 s 567884 -800 567996 480 0 la_oenb[124]
port 447 nsew signal input
rlabel metal2 s 571430 -800 571542 480 0 la_oenb[125]
port 448 nsew signal input
rlabel metal2 s 574976 -800 575088 480 0 la_oenb[126]
port 449 nsew signal input
rlabel metal2 s 578522 -800 578634 480 0 la_oenb[127]
port 450 nsew signal input
rlabel metal2 s 170732 -800 170844 480 0 la_oenb[12]
port 451 nsew signal input
rlabel metal2 s 174278 -800 174390 480 0 la_oenb[13]
port 452 nsew signal input
rlabel metal2 s 177824 -800 177936 480 0 la_oenb[14]
port 453 nsew signal input
rlabel metal2 s 181370 -800 181482 480 0 la_oenb[15]
port 454 nsew signal input
rlabel metal2 s 184916 -800 185028 480 0 la_oenb[16]
port 455 nsew signal input
rlabel metal2 s 188462 -800 188574 480 0 la_oenb[17]
port 456 nsew signal input
rlabel metal2 s 192008 -800 192120 480 0 la_oenb[18]
port 457 nsew signal input
rlabel metal2 s 195554 -800 195666 480 0 la_oenb[19]
port 458 nsew signal input
rlabel metal2 s 131726 -800 131838 480 0 la_oenb[1]
port 459 nsew signal input
rlabel metal2 s 199100 -800 199212 480 0 la_oenb[20]
port 460 nsew signal input
rlabel metal2 s 202646 -800 202758 480 0 la_oenb[21]
port 461 nsew signal input
rlabel metal2 s 206192 -800 206304 480 0 la_oenb[22]
port 462 nsew signal input
rlabel metal2 s 209738 -800 209850 480 0 la_oenb[23]
port 463 nsew signal input
rlabel metal2 s 213284 -800 213396 480 0 la_oenb[24]
port 464 nsew signal input
rlabel metal2 s 216830 -800 216942 480 0 la_oenb[25]
port 465 nsew signal input
rlabel metal2 s 220376 -800 220488 480 0 la_oenb[26]
port 466 nsew signal input
rlabel metal2 s 223922 -800 224034 480 0 la_oenb[27]
port 467 nsew signal input
rlabel metal2 s 227468 -800 227580 480 0 la_oenb[28]
port 468 nsew signal input
rlabel metal2 s 231014 -800 231126 480 0 la_oenb[29]
port 469 nsew signal input
rlabel metal2 s 135272 -800 135384 480 0 la_oenb[2]
port 470 nsew signal input
rlabel metal2 s 234560 -800 234672 480 0 la_oenb[30]
port 471 nsew signal input
rlabel metal2 s 238106 -800 238218 480 0 la_oenb[31]
port 472 nsew signal input
rlabel metal2 s 241652 -800 241764 480 0 la_oenb[32]
port 473 nsew signal input
rlabel metal2 s 245198 -800 245310 480 0 la_oenb[33]
port 474 nsew signal input
rlabel metal2 s 248744 -800 248856 480 0 la_oenb[34]
port 475 nsew signal input
rlabel metal2 s 252290 -800 252402 480 0 la_oenb[35]
port 476 nsew signal input
rlabel metal2 s 255836 -800 255948 480 0 la_oenb[36]
port 477 nsew signal input
rlabel metal2 s 259382 -800 259494 480 0 la_oenb[37]
port 478 nsew signal input
rlabel metal2 s 262928 -800 263040 480 0 la_oenb[38]
port 479 nsew signal input
rlabel metal2 s 266474 -800 266586 480 0 la_oenb[39]
port 480 nsew signal input
rlabel metal2 s 138818 -800 138930 480 0 la_oenb[3]
port 481 nsew signal input
rlabel metal2 s 270020 -800 270132 480 0 la_oenb[40]
port 482 nsew signal input
rlabel metal2 s 273566 -800 273678 480 0 la_oenb[41]
port 483 nsew signal input
rlabel metal2 s 277112 -800 277224 480 0 la_oenb[42]
port 484 nsew signal input
rlabel metal2 s 280658 -800 280770 480 0 la_oenb[43]
port 485 nsew signal input
rlabel metal2 s 284204 -800 284316 480 0 la_oenb[44]
port 486 nsew signal input
rlabel metal2 s 287750 -800 287862 480 0 la_oenb[45]
port 487 nsew signal input
rlabel metal2 s 291296 -800 291408 480 0 la_oenb[46]
port 488 nsew signal input
rlabel metal2 s 294842 -800 294954 480 0 la_oenb[47]
port 489 nsew signal input
rlabel metal2 s 298388 -800 298500 480 0 la_oenb[48]
port 490 nsew signal input
rlabel metal2 s 301934 -800 302046 480 0 la_oenb[49]
port 491 nsew signal input
rlabel metal2 s 142364 -800 142476 480 0 la_oenb[4]
port 492 nsew signal input
rlabel metal2 s 305480 -800 305592 480 0 la_oenb[50]
port 493 nsew signal input
rlabel metal2 s 309026 -800 309138 480 0 la_oenb[51]
port 494 nsew signal input
rlabel metal2 s 312572 -800 312684 480 0 la_oenb[52]
port 495 nsew signal input
rlabel metal2 s 316118 -800 316230 480 0 la_oenb[53]
port 496 nsew signal input
rlabel metal2 s 319664 -800 319776 480 0 la_oenb[54]
port 497 nsew signal input
rlabel metal2 s 323210 -800 323322 480 0 la_oenb[55]
port 498 nsew signal input
rlabel metal2 s 326756 -800 326868 480 0 la_oenb[56]
port 499 nsew signal input
rlabel metal2 s 330302 -800 330414 480 0 la_oenb[57]
port 500 nsew signal input
rlabel metal2 s 333848 -800 333960 480 0 la_oenb[58]
port 501 nsew signal input
rlabel metal2 s 337394 -800 337506 480 0 la_oenb[59]
port 502 nsew signal input
rlabel metal2 s 145910 -800 146022 480 0 la_oenb[5]
port 503 nsew signal input
rlabel metal2 s 340940 -800 341052 480 0 la_oenb[60]
port 504 nsew signal input
rlabel metal2 s 344486 -800 344598 480 0 la_oenb[61]
port 505 nsew signal input
rlabel metal2 s 348032 -800 348144 480 0 la_oenb[62]
port 506 nsew signal input
rlabel metal2 s 351578 -800 351690 480 0 la_oenb[63]
port 507 nsew signal input
rlabel metal2 s 355124 -800 355236 480 0 la_oenb[64]
port 508 nsew signal input
rlabel metal2 s 358670 -800 358782 480 0 la_oenb[65]
port 509 nsew signal input
rlabel metal2 s 362216 -800 362328 480 0 la_oenb[66]
port 510 nsew signal input
rlabel metal2 s 365762 -800 365874 480 0 la_oenb[67]
port 511 nsew signal input
rlabel metal2 s 369308 -800 369420 480 0 la_oenb[68]
port 512 nsew signal input
rlabel metal2 s 372854 -800 372966 480 0 la_oenb[69]
port 513 nsew signal input
rlabel metal2 s 149456 -800 149568 480 0 la_oenb[6]
port 514 nsew signal input
rlabel metal2 s 376400 -800 376512 480 0 la_oenb[70]
port 515 nsew signal input
rlabel metal2 s 379946 -800 380058 480 0 la_oenb[71]
port 516 nsew signal input
rlabel metal2 s 383492 -800 383604 480 0 la_oenb[72]
port 517 nsew signal input
rlabel metal2 s 387038 -800 387150 480 0 la_oenb[73]
port 518 nsew signal input
rlabel metal2 s 390584 -800 390696 480 0 la_oenb[74]
port 519 nsew signal input
rlabel metal2 s 394130 -800 394242 480 0 la_oenb[75]
port 520 nsew signal input
rlabel metal2 s 397676 -800 397788 480 0 la_oenb[76]
port 521 nsew signal input
rlabel metal2 s 401222 -800 401334 480 0 la_oenb[77]
port 522 nsew signal input
rlabel metal2 s 404768 -800 404880 480 0 la_oenb[78]
port 523 nsew signal input
rlabel metal2 s 408314 -800 408426 480 0 la_oenb[79]
port 524 nsew signal input
rlabel metal2 s 153002 -800 153114 480 0 la_oenb[7]
port 525 nsew signal input
rlabel metal2 s 411860 -800 411972 480 0 la_oenb[80]
port 526 nsew signal input
rlabel metal2 s 415406 -800 415518 480 0 la_oenb[81]
port 527 nsew signal input
rlabel metal2 s 418952 -800 419064 480 0 la_oenb[82]
port 528 nsew signal input
rlabel metal2 s 422498 -800 422610 480 0 la_oenb[83]
port 529 nsew signal input
rlabel metal2 s 426044 -800 426156 480 0 la_oenb[84]
port 530 nsew signal input
rlabel metal2 s 429590 -800 429702 480 0 la_oenb[85]
port 531 nsew signal input
rlabel metal2 s 433136 -800 433248 480 0 la_oenb[86]
port 532 nsew signal input
rlabel metal2 s 436682 -800 436794 480 0 la_oenb[87]
port 533 nsew signal input
rlabel metal2 s 440228 -800 440340 480 0 la_oenb[88]
port 534 nsew signal input
rlabel metal2 s 443774 -800 443886 480 0 la_oenb[89]
port 535 nsew signal input
rlabel metal2 s 156548 -800 156660 480 0 la_oenb[8]
port 536 nsew signal input
rlabel metal2 s 447320 -800 447432 480 0 la_oenb[90]
port 537 nsew signal input
rlabel metal2 s 450866 -800 450978 480 0 la_oenb[91]
port 538 nsew signal input
rlabel metal2 s 454412 -800 454524 480 0 la_oenb[92]
port 539 nsew signal input
rlabel metal2 s 457958 -800 458070 480 0 la_oenb[93]
port 540 nsew signal input
rlabel metal2 s 461504 -800 461616 480 0 la_oenb[94]
port 541 nsew signal input
rlabel metal2 s 465050 -800 465162 480 0 la_oenb[95]
port 542 nsew signal input
rlabel metal2 s 468596 -800 468708 480 0 la_oenb[96]
port 543 nsew signal input
rlabel metal2 s 472142 -800 472254 480 0 la_oenb[97]
port 544 nsew signal input
rlabel metal2 s 475688 -800 475800 480 0 la_oenb[98]
port 545 nsew signal input
rlabel metal2 s 479234 -800 479346 480 0 la_oenb[99]
port 546 nsew signal input
rlabel metal2 s 160094 -800 160206 480 0 la_oenb[9]
port 547 nsew signal input
rlabel metal2 s 579704 -800 579816 480 0 user_clock2
port 548 nsew signal input
rlabel metal2 s 580886 -800 580998 480 0 user_irq[0]
port 549 nsew signal tristate
rlabel metal2 s 582068 -800 582180 480 0 user_irq[1]
port 550 nsew signal tristate
rlabel metal2 s 583250 -800 583362 480 0 user_irq[2]
port 551 nsew signal tristate
rlabel metal3 s 582340 639784 584800 644584 0 vccd1
port 552 nsew signal bidirectional
rlabel metal3 s 582340 629784 584800 634584 0 vccd1
port 553 nsew signal bidirectional
rlabel metal3 s 0 643842 1660 648642 0 vccd2
port 554 nsew signal bidirectional
rlabel metal3 s 0 633842 1660 638642 0 vccd2
port 555 nsew signal bidirectional
rlabel metal3 s 582340 540562 584800 545362 0 vdda1
port 556 nsew signal bidirectional
rlabel metal3 s 582340 550562 584800 555362 0 vdda1
port 557 nsew signal bidirectional
rlabel metal3 s 582340 235230 584800 240030 0 vdda1
port 558 nsew signal bidirectional
rlabel metal3 s 582340 225230 584800 230030 0 vdda1
port 559 nsew signal bidirectional
rlabel metal3 s 0 204888 1660 209688 0 vdda2
port 560 nsew signal bidirectional
rlabel metal3 s 0 214888 1660 219688 0 vdda2
port 561 nsew signal bidirectional
rlabel metal3 s 520594 702340 525394 704800 0 vssa1
port 562 nsew signal bidirectional
rlabel metal3 s 510594 702340 515394 704800 0 vssa1
port 563 nsew signal bidirectional
rlabel metal3 s 582340 146830 584800 151630 0 vssa1
port 564 nsew signal bidirectional
rlabel metal3 s 582340 136830 584800 141630 0 vssa1
port 565 nsew signal bidirectional
rlabel metal3 s 0 559442 1660 564242 0 vssa2
port 566 nsew signal bidirectional
rlabel metal3 s 0 549442 1660 554242 0 vssa2
port 567 nsew signal bidirectional
rlabel metal3 s 582340 191430 584800 196230 0 vssd1
port 568 nsew signal bidirectional
rlabel metal3 s 582340 181430 584800 186230 0 vssd1
port 569 nsew signal bidirectional
rlabel metal3 s 0 172888 1660 177688 0 vssd2
port 570 nsew signal bidirectional
rlabel metal3 s 0 162888 1660 167688 0 vssd2
port 571 nsew signal bidirectional
rlabel metal2 s 524 -800 636 480 0 wb_clk_i
port 572 nsew signal input
rlabel metal2 s 1706 -800 1818 480 0 wb_rst_i
port 573 nsew signal input
rlabel metal2 s 2888 -800 3000 480 0 wbs_ack_o
port 574 nsew signal tristate
rlabel metal2 s 7616 -800 7728 480 0 wbs_adr_i[0]
port 575 nsew signal input
rlabel metal2 s 47804 -800 47916 480 0 wbs_adr_i[10]
port 576 nsew signal input
rlabel metal2 s 51350 -800 51462 480 0 wbs_adr_i[11]
port 577 nsew signal input
rlabel metal2 s 54896 -800 55008 480 0 wbs_adr_i[12]
port 578 nsew signal input
rlabel metal2 s 58442 -800 58554 480 0 wbs_adr_i[13]
port 579 nsew signal input
rlabel metal2 s 61988 -800 62100 480 0 wbs_adr_i[14]
port 580 nsew signal input
rlabel metal2 s 65534 -800 65646 480 0 wbs_adr_i[15]
port 581 nsew signal input
rlabel metal2 s 69080 -800 69192 480 0 wbs_adr_i[16]
port 582 nsew signal input
rlabel metal2 s 72626 -800 72738 480 0 wbs_adr_i[17]
port 583 nsew signal input
rlabel metal2 s 76172 -800 76284 480 0 wbs_adr_i[18]
port 584 nsew signal input
rlabel metal2 s 79718 -800 79830 480 0 wbs_adr_i[19]
port 585 nsew signal input
rlabel metal2 s 12344 -800 12456 480 0 wbs_adr_i[1]
port 586 nsew signal input
rlabel metal2 s 83264 -800 83376 480 0 wbs_adr_i[20]
port 587 nsew signal input
rlabel metal2 s 86810 -800 86922 480 0 wbs_adr_i[21]
port 588 nsew signal input
rlabel metal2 s 90356 -800 90468 480 0 wbs_adr_i[22]
port 589 nsew signal input
rlabel metal2 s 93902 -800 94014 480 0 wbs_adr_i[23]
port 590 nsew signal input
rlabel metal2 s 97448 -800 97560 480 0 wbs_adr_i[24]
port 591 nsew signal input
rlabel metal2 s 100994 -800 101106 480 0 wbs_adr_i[25]
port 592 nsew signal input
rlabel metal2 s 104540 -800 104652 480 0 wbs_adr_i[26]
port 593 nsew signal input
rlabel metal2 s 108086 -800 108198 480 0 wbs_adr_i[27]
port 594 nsew signal input
rlabel metal2 s 111632 -800 111744 480 0 wbs_adr_i[28]
port 595 nsew signal input
rlabel metal2 s 115178 -800 115290 480 0 wbs_adr_i[29]
port 596 nsew signal input
rlabel metal2 s 17072 -800 17184 480 0 wbs_adr_i[2]
port 597 nsew signal input
rlabel metal2 s 118724 -800 118836 480 0 wbs_adr_i[30]
port 598 nsew signal input
rlabel metal2 s 122270 -800 122382 480 0 wbs_adr_i[31]
port 599 nsew signal input
rlabel metal2 s 21800 -800 21912 480 0 wbs_adr_i[3]
port 600 nsew signal input
rlabel metal2 s 26528 -800 26640 480 0 wbs_adr_i[4]
port 601 nsew signal input
rlabel metal2 s 30074 -800 30186 480 0 wbs_adr_i[5]
port 602 nsew signal input
rlabel metal2 s 33620 -800 33732 480 0 wbs_adr_i[6]
port 603 nsew signal input
rlabel metal2 s 37166 -800 37278 480 0 wbs_adr_i[7]
port 604 nsew signal input
rlabel metal2 s 40712 -800 40824 480 0 wbs_adr_i[8]
port 605 nsew signal input
rlabel metal2 s 44258 -800 44370 480 0 wbs_adr_i[9]
port 606 nsew signal input
rlabel metal2 s 4070 -800 4182 480 0 wbs_cyc_i
port 607 nsew signal input
rlabel metal2 s 8798 -800 8910 480 0 wbs_dat_i[0]
port 608 nsew signal input
rlabel metal2 s 48986 -800 49098 480 0 wbs_dat_i[10]
port 609 nsew signal input
rlabel metal2 s 52532 -800 52644 480 0 wbs_dat_i[11]
port 610 nsew signal input
rlabel metal2 s 56078 -800 56190 480 0 wbs_dat_i[12]
port 611 nsew signal input
rlabel metal2 s 59624 -800 59736 480 0 wbs_dat_i[13]
port 612 nsew signal input
rlabel metal2 s 63170 -800 63282 480 0 wbs_dat_i[14]
port 613 nsew signal input
rlabel metal2 s 66716 -800 66828 480 0 wbs_dat_i[15]
port 614 nsew signal input
rlabel metal2 s 70262 -800 70374 480 0 wbs_dat_i[16]
port 615 nsew signal input
rlabel metal2 s 73808 -800 73920 480 0 wbs_dat_i[17]
port 616 nsew signal input
rlabel metal2 s 77354 -800 77466 480 0 wbs_dat_i[18]
port 617 nsew signal input
rlabel metal2 s 80900 -800 81012 480 0 wbs_dat_i[19]
port 618 nsew signal input
rlabel metal2 s 13526 -800 13638 480 0 wbs_dat_i[1]
port 619 nsew signal input
rlabel metal2 s 84446 -800 84558 480 0 wbs_dat_i[20]
port 620 nsew signal input
rlabel metal2 s 87992 -800 88104 480 0 wbs_dat_i[21]
port 621 nsew signal input
rlabel metal2 s 91538 -800 91650 480 0 wbs_dat_i[22]
port 622 nsew signal input
rlabel metal2 s 95084 -800 95196 480 0 wbs_dat_i[23]
port 623 nsew signal input
rlabel metal2 s 98630 -800 98742 480 0 wbs_dat_i[24]
port 624 nsew signal input
rlabel metal2 s 102176 -800 102288 480 0 wbs_dat_i[25]
port 625 nsew signal input
rlabel metal2 s 105722 -800 105834 480 0 wbs_dat_i[26]
port 626 nsew signal input
rlabel metal2 s 109268 -800 109380 480 0 wbs_dat_i[27]
port 627 nsew signal input
rlabel metal2 s 112814 -800 112926 480 0 wbs_dat_i[28]
port 628 nsew signal input
rlabel metal2 s 116360 -800 116472 480 0 wbs_dat_i[29]
port 629 nsew signal input
rlabel metal2 s 18254 -800 18366 480 0 wbs_dat_i[2]
port 630 nsew signal input
rlabel metal2 s 119906 -800 120018 480 0 wbs_dat_i[30]
port 631 nsew signal input
rlabel metal2 s 123452 -800 123564 480 0 wbs_dat_i[31]
port 632 nsew signal input
rlabel metal2 s 22982 -800 23094 480 0 wbs_dat_i[3]
port 633 nsew signal input
rlabel metal2 s 27710 -800 27822 480 0 wbs_dat_i[4]
port 634 nsew signal input
rlabel metal2 s 31256 -800 31368 480 0 wbs_dat_i[5]
port 635 nsew signal input
rlabel metal2 s 34802 -800 34914 480 0 wbs_dat_i[6]
port 636 nsew signal input
rlabel metal2 s 38348 -800 38460 480 0 wbs_dat_i[7]
port 637 nsew signal input
rlabel metal2 s 41894 -800 42006 480 0 wbs_dat_i[8]
port 638 nsew signal input
rlabel metal2 s 45440 -800 45552 480 0 wbs_dat_i[9]
port 639 nsew signal input
rlabel metal2 s 9980 -800 10092 480 0 wbs_dat_o[0]
port 640 nsew signal tristate
rlabel metal2 s 50168 -800 50280 480 0 wbs_dat_o[10]
port 641 nsew signal tristate
rlabel metal2 s 53714 -800 53826 480 0 wbs_dat_o[11]
port 642 nsew signal tristate
rlabel metal2 s 57260 -800 57372 480 0 wbs_dat_o[12]
port 643 nsew signal tristate
rlabel metal2 s 60806 -800 60918 480 0 wbs_dat_o[13]
port 644 nsew signal tristate
rlabel metal2 s 64352 -800 64464 480 0 wbs_dat_o[14]
port 645 nsew signal tristate
rlabel metal2 s 67898 -800 68010 480 0 wbs_dat_o[15]
port 646 nsew signal tristate
rlabel metal2 s 71444 -800 71556 480 0 wbs_dat_o[16]
port 647 nsew signal tristate
rlabel metal2 s 74990 -800 75102 480 0 wbs_dat_o[17]
port 648 nsew signal tristate
rlabel metal2 s 78536 -800 78648 480 0 wbs_dat_o[18]
port 649 nsew signal tristate
rlabel metal2 s 82082 -800 82194 480 0 wbs_dat_o[19]
port 650 nsew signal tristate
rlabel metal2 s 14708 -800 14820 480 0 wbs_dat_o[1]
port 651 nsew signal tristate
rlabel metal2 s 85628 -800 85740 480 0 wbs_dat_o[20]
port 652 nsew signal tristate
rlabel metal2 s 89174 -800 89286 480 0 wbs_dat_o[21]
port 653 nsew signal tristate
rlabel metal2 s 92720 -800 92832 480 0 wbs_dat_o[22]
port 654 nsew signal tristate
rlabel metal2 s 96266 -800 96378 480 0 wbs_dat_o[23]
port 655 nsew signal tristate
rlabel metal2 s 99812 -800 99924 480 0 wbs_dat_o[24]
port 656 nsew signal tristate
rlabel metal2 s 103358 -800 103470 480 0 wbs_dat_o[25]
port 657 nsew signal tristate
rlabel metal2 s 106904 -800 107016 480 0 wbs_dat_o[26]
port 658 nsew signal tristate
rlabel metal2 s 110450 -800 110562 480 0 wbs_dat_o[27]
port 659 nsew signal tristate
rlabel metal2 s 113996 -800 114108 480 0 wbs_dat_o[28]
port 660 nsew signal tristate
rlabel metal2 s 117542 -800 117654 480 0 wbs_dat_o[29]
port 661 nsew signal tristate
rlabel metal2 s 19436 -800 19548 480 0 wbs_dat_o[2]
port 662 nsew signal tristate
rlabel metal2 s 121088 -800 121200 480 0 wbs_dat_o[30]
port 663 nsew signal tristate
rlabel metal2 s 124634 -800 124746 480 0 wbs_dat_o[31]
port 664 nsew signal tristate
rlabel metal2 s 24164 -800 24276 480 0 wbs_dat_o[3]
port 665 nsew signal tristate
rlabel metal2 s 28892 -800 29004 480 0 wbs_dat_o[4]
port 666 nsew signal tristate
rlabel metal2 s 32438 -800 32550 480 0 wbs_dat_o[5]
port 667 nsew signal tristate
rlabel metal2 s 35984 -800 36096 480 0 wbs_dat_o[6]
port 668 nsew signal tristate
rlabel metal2 s 39530 -800 39642 480 0 wbs_dat_o[7]
port 669 nsew signal tristate
rlabel metal2 s 43076 -800 43188 480 0 wbs_dat_o[8]
port 670 nsew signal tristate
rlabel metal2 s 46622 -800 46734 480 0 wbs_dat_o[9]
port 671 nsew signal tristate
rlabel metal2 s 11162 -800 11274 480 0 wbs_sel_i[0]
port 672 nsew signal input
rlabel metal2 s 15890 -800 16002 480 0 wbs_sel_i[1]
port 673 nsew signal input
rlabel metal2 s 20618 -800 20730 480 0 wbs_sel_i[2]
port 674 nsew signal input
rlabel metal2 s 25346 -800 25458 480 0 wbs_sel_i[3]
port 675 nsew signal input
rlabel metal2 s 5252 -800 5364 480 0 wbs_stb_i
port 676 nsew signal input
rlabel metal2 s 6434 -800 6546 480 0 wbs_we_i
port 677 nsew signal input
rlabel space 26080 559400 65590 564330 0 GND
rlabel metal2 56720 466080 56860 660460 1 CTRL2
rlabel metal2 56480 421660 56620 660980 1 CTRL3
rlabel metal2 56200 378460 56340 661580 1 CTRL4
rlabel metal1 14920 668060 15420 682040 0 VCTRL
rlabel metal3 17070 688210 41870 689330 1 OUT0
rlabel metal3 43180 688360 70760 689480 1 OUT180
rlabel metal3 163400 360000 198200 362000 0 txinb
rlabel metal3 163400 466000 198200 468000 0 txina
rlabel metal2 56980 508120 57120 660100 1 CTRL1
rlabel metal4 22200 605800 23800 611800 0 REF
rlabel metal2 55960 335420 56100 662700 1 CTRL5
rlabel metal2 148200 430920 148420 435520 0 REF2
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
