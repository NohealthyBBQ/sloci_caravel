magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -1887 181 -1825 187
rect -1759 181 -1697 187
rect -1631 181 -1569 187
rect -1503 181 -1441 187
rect -1375 181 -1313 187
rect -1247 181 -1185 187
rect -1119 181 -1057 187
rect -991 181 -929 187
rect -863 181 -801 187
rect -735 181 -673 187
rect -607 181 -545 187
rect -479 181 -417 187
rect -351 181 -289 187
rect -223 181 -161 187
rect -95 181 -33 187
rect 33 181 95 187
rect 161 181 223 187
rect 289 181 351 187
rect 417 181 479 187
rect 545 181 607 187
rect 673 181 735 187
rect 801 181 863 187
rect 929 181 991 187
rect 1057 181 1119 187
rect 1185 181 1247 187
rect 1313 181 1375 187
rect 1441 181 1503 187
rect 1569 181 1631 187
rect 1697 181 1759 187
rect 1825 181 1887 187
rect -1887 147 -1873 181
rect -1759 147 -1745 181
rect -1631 147 -1617 181
rect -1503 147 -1489 181
rect -1375 147 -1361 181
rect -1247 147 -1233 181
rect -1119 147 -1105 181
rect -991 147 -977 181
rect -863 147 -849 181
rect -735 147 -721 181
rect -607 147 -593 181
rect -479 147 -465 181
rect -351 147 -337 181
rect -223 147 -209 181
rect -95 147 -81 181
rect 33 147 47 181
rect 161 147 175 181
rect 289 147 303 181
rect 417 147 431 181
rect 545 147 559 181
rect 673 147 687 181
rect 801 147 815 181
rect 929 147 943 181
rect 1057 147 1071 181
rect 1185 147 1199 181
rect 1313 147 1327 181
rect 1441 147 1455 181
rect 1569 147 1583 181
rect 1697 147 1711 181
rect 1825 147 1839 181
rect -1887 141 -1825 147
rect -1759 141 -1697 147
rect -1631 141 -1569 147
rect -1503 141 -1441 147
rect -1375 141 -1313 147
rect -1247 141 -1185 147
rect -1119 141 -1057 147
rect -991 141 -929 147
rect -863 141 -801 147
rect -735 141 -673 147
rect -607 141 -545 147
rect -479 141 -417 147
rect -351 141 -289 147
rect -223 141 -161 147
rect -95 141 -33 147
rect 33 141 95 147
rect 161 141 223 147
rect 289 141 351 147
rect 417 141 479 147
rect 545 141 607 147
rect 673 141 735 147
rect 801 141 863 147
rect 929 141 991 147
rect 1057 141 1119 147
rect 1185 141 1247 147
rect 1313 141 1375 147
rect 1441 141 1503 147
rect 1569 141 1631 147
rect 1697 141 1759 147
rect 1825 141 1887 147
rect -1887 -147 -1825 -141
rect -1759 -147 -1697 -141
rect -1631 -147 -1569 -141
rect -1503 -147 -1441 -141
rect -1375 -147 -1313 -141
rect -1247 -147 -1185 -141
rect -1119 -147 -1057 -141
rect -991 -147 -929 -141
rect -863 -147 -801 -141
rect -735 -147 -673 -141
rect -607 -147 -545 -141
rect -479 -147 -417 -141
rect -351 -147 -289 -141
rect -223 -147 -161 -141
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect 161 -147 223 -141
rect 289 -147 351 -141
rect 417 -147 479 -141
rect 545 -147 607 -141
rect 673 -147 735 -141
rect 801 -147 863 -141
rect 929 -147 991 -141
rect 1057 -147 1119 -141
rect 1185 -147 1247 -141
rect 1313 -147 1375 -141
rect 1441 -147 1503 -141
rect 1569 -147 1631 -141
rect 1697 -147 1759 -141
rect 1825 -147 1887 -141
rect -1887 -181 -1873 -147
rect -1759 -181 -1745 -147
rect -1631 -181 -1617 -147
rect -1503 -181 -1489 -147
rect -1375 -181 -1361 -147
rect -1247 -181 -1233 -147
rect -1119 -181 -1105 -147
rect -991 -181 -977 -147
rect -863 -181 -849 -147
rect -735 -181 -721 -147
rect -607 -181 -593 -147
rect -479 -181 -465 -147
rect -351 -181 -337 -147
rect -223 -181 -209 -147
rect -95 -181 -81 -147
rect 33 -181 47 -147
rect 161 -181 175 -147
rect 289 -181 303 -147
rect 417 -181 431 -147
rect 545 -181 559 -147
rect 673 -181 687 -147
rect 801 -181 815 -147
rect 929 -181 943 -147
rect 1057 -181 1071 -147
rect 1185 -181 1199 -147
rect 1313 -181 1327 -147
rect 1441 -181 1455 -147
rect 1569 -181 1583 -147
rect 1697 -181 1711 -147
rect 1825 -181 1839 -147
rect -1887 -187 -1825 -181
rect -1759 -187 -1697 -181
rect -1631 -187 -1569 -181
rect -1503 -187 -1441 -181
rect -1375 -187 -1313 -181
rect -1247 -187 -1185 -181
rect -1119 -187 -1057 -181
rect -991 -187 -929 -181
rect -863 -187 -801 -181
rect -735 -187 -673 -181
rect -607 -187 -545 -181
rect -479 -187 -417 -181
rect -351 -187 -289 -181
rect -223 -187 -161 -181
rect -95 -187 -33 -181
rect 33 -187 95 -181
rect 161 -187 223 -181
rect 289 -187 351 -181
rect 417 -187 479 -181
rect 545 -187 607 -181
rect 673 -187 735 -181
rect 801 -187 863 -181
rect 929 -187 991 -181
rect 1057 -187 1119 -181
rect 1185 -187 1247 -181
rect 1313 -187 1375 -181
rect 1441 -187 1503 -181
rect 1569 -187 1631 -181
rect 1697 -187 1759 -181
rect 1825 -187 1887 -181
<< nwell >>
rect -2087 -319 2087 319
<< pmoslvt >>
rect -1891 -100 -1821 100
rect -1763 -100 -1693 100
rect -1635 -100 -1565 100
rect -1507 -100 -1437 100
rect -1379 -100 -1309 100
rect -1251 -100 -1181 100
rect -1123 -100 -1053 100
rect -995 -100 -925 100
rect -867 -100 -797 100
rect -739 -100 -669 100
rect -611 -100 -541 100
rect -483 -100 -413 100
rect -355 -100 -285 100
rect -227 -100 -157 100
rect -99 -100 -29 100
rect 29 -100 99 100
rect 157 -100 227 100
rect 285 -100 355 100
rect 413 -100 483 100
rect 541 -100 611 100
rect 669 -100 739 100
rect 797 -100 867 100
rect 925 -100 995 100
rect 1053 -100 1123 100
rect 1181 -100 1251 100
rect 1309 -100 1379 100
rect 1437 -100 1507 100
rect 1565 -100 1635 100
rect 1693 -100 1763 100
rect 1821 -100 1891 100
<< pdiff >>
rect -1949 85 -1891 100
rect -1949 51 -1937 85
rect -1903 51 -1891 85
rect -1949 17 -1891 51
rect -1949 -17 -1937 17
rect -1903 -17 -1891 17
rect -1949 -51 -1891 -17
rect -1949 -85 -1937 -51
rect -1903 -85 -1891 -51
rect -1949 -100 -1891 -85
rect -1821 85 -1763 100
rect -1821 51 -1809 85
rect -1775 51 -1763 85
rect -1821 17 -1763 51
rect -1821 -17 -1809 17
rect -1775 -17 -1763 17
rect -1821 -51 -1763 -17
rect -1821 -85 -1809 -51
rect -1775 -85 -1763 -51
rect -1821 -100 -1763 -85
rect -1693 85 -1635 100
rect -1693 51 -1681 85
rect -1647 51 -1635 85
rect -1693 17 -1635 51
rect -1693 -17 -1681 17
rect -1647 -17 -1635 17
rect -1693 -51 -1635 -17
rect -1693 -85 -1681 -51
rect -1647 -85 -1635 -51
rect -1693 -100 -1635 -85
rect -1565 85 -1507 100
rect -1565 51 -1553 85
rect -1519 51 -1507 85
rect -1565 17 -1507 51
rect -1565 -17 -1553 17
rect -1519 -17 -1507 17
rect -1565 -51 -1507 -17
rect -1565 -85 -1553 -51
rect -1519 -85 -1507 -51
rect -1565 -100 -1507 -85
rect -1437 85 -1379 100
rect -1437 51 -1425 85
rect -1391 51 -1379 85
rect -1437 17 -1379 51
rect -1437 -17 -1425 17
rect -1391 -17 -1379 17
rect -1437 -51 -1379 -17
rect -1437 -85 -1425 -51
rect -1391 -85 -1379 -51
rect -1437 -100 -1379 -85
rect -1309 85 -1251 100
rect -1309 51 -1297 85
rect -1263 51 -1251 85
rect -1309 17 -1251 51
rect -1309 -17 -1297 17
rect -1263 -17 -1251 17
rect -1309 -51 -1251 -17
rect -1309 -85 -1297 -51
rect -1263 -85 -1251 -51
rect -1309 -100 -1251 -85
rect -1181 85 -1123 100
rect -1181 51 -1169 85
rect -1135 51 -1123 85
rect -1181 17 -1123 51
rect -1181 -17 -1169 17
rect -1135 -17 -1123 17
rect -1181 -51 -1123 -17
rect -1181 -85 -1169 -51
rect -1135 -85 -1123 -51
rect -1181 -100 -1123 -85
rect -1053 85 -995 100
rect -1053 51 -1041 85
rect -1007 51 -995 85
rect -1053 17 -995 51
rect -1053 -17 -1041 17
rect -1007 -17 -995 17
rect -1053 -51 -995 -17
rect -1053 -85 -1041 -51
rect -1007 -85 -995 -51
rect -1053 -100 -995 -85
rect -925 85 -867 100
rect -925 51 -913 85
rect -879 51 -867 85
rect -925 17 -867 51
rect -925 -17 -913 17
rect -879 -17 -867 17
rect -925 -51 -867 -17
rect -925 -85 -913 -51
rect -879 -85 -867 -51
rect -925 -100 -867 -85
rect -797 85 -739 100
rect -797 51 -785 85
rect -751 51 -739 85
rect -797 17 -739 51
rect -797 -17 -785 17
rect -751 -17 -739 17
rect -797 -51 -739 -17
rect -797 -85 -785 -51
rect -751 -85 -739 -51
rect -797 -100 -739 -85
rect -669 85 -611 100
rect -669 51 -657 85
rect -623 51 -611 85
rect -669 17 -611 51
rect -669 -17 -657 17
rect -623 -17 -611 17
rect -669 -51 -611 -17
rect -669 -85 -657 -51
rect -623 -85 -611 -51
rect -669 -100 -611 -85
rect -541 85 -483 100
rect -541 51 -529 85
rect -495 51 -483 85
rect -541 17 -483 51
rect -541 -17 -529 17
rect -495 -17 -483 17
rect -541 -51 -483 -17
rect -541 -85 -529 -51
rect -495 -85 -483 -51
rect -541 -100 -483 -85
rect -413 85 -355 100
rect -413 51 -401 85
rect -367 51 -355 85
rect -413 17 -355 51
rect -413 -17 -401 17
rect -367 -17 -355 17
rect -413 -51 -355 -17
rect -413 -85 -401 -51
rect -367 -85 -355 -51
rect -413 -100 -355 -85
rect -285 85 -227 100
rect -285 51 -273 85
rect -239 51 -227 85
rect -285 17 -227 51
rect -285 -17 -273 17
rect -239 -17 -227 17
rect -285 -51 -227 -17
rect -285 -85 -273 -51
rect -239 -85 -227 -51
rect -285 -100 -227 -85
rect -157 85 -99 100
rect -157 51 -145 85
rect -111 51 -99 85
rect -157 17 -99 51
rect -157 -17 -145 17
rect -111 -17 -99 17
rect -157 -51 -99 -17
rect -157 -85 -145 -51
rect -111 -85 -99 -51
rect -157 -100 -99 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 99 85 157 100
rect 99 51 111 85
rect 145 51 157 85
rect 99 17 157 51
rect 99 -17 111 17
rect 145 -17 157 17
rect 99 -51 157 -17
rect 99 -85 111 -51
rect 145 -85 157 -51
rect 99 -100 157 -85
rect 227 85 285 100
rect 227 51 239 85
rect 273 51 285 85
rect 227 17 285 51
rect 227 -17 239 17
rect 273 -17 285 17
rect 227 -51 285 -17
rect 227 -85 239 -51
rect 273 -85 285 -51
rect 227 -100 285 -85
rect 355 85 413 100
rect 355 51 367 85
rect 401 51 413 85
rect 355 17 413 51
rect 355 -17 367 17
rect 401 -17 413 17
rect 355 -51 413 -17
rect 355 -85 367 -51
rect 401 -85 413 -51
rect 355 -100 413 -85
rect 483 85 541 100
rect 483 51 495 85
rect 529 51 541 85
rect 483 17 541 51
rect 483 -17 495 17
rect 529 -17 541 17
rect 483 -51 541 -17
rect 483 -85 495 -51
rect 529 -85 541 -51
rect 483 -100 541 -85
rect 611 85 669 100
rect 611 51 623 85
rect 657 51 669 85
rect 611 17 669 51
rect 611 -17 623 17
rect 657 -17 669 17
rect 611 -51 669 -17
rect 611 -85 623 -51
rect 657 -85 669 -51
rect 611 -100 669 -85
rect 739 85 797 100
rect 739 51 751 85
rect 785 51 797 85
rect 739 17 797 51
rect 739 -17 751 17
rect 785 -17 797 17
rect 739 -51 797 -17
rect 739 -85 751 -51
rect 785 -85 797 -51
rect 739 -100 797 -85
rect 867 85 925 100
rect 867 51 879 85
rect 913 51 925 85
rect 867 17 925 51
rect 867 -17 879 17
rect 913 -17 925 17
rect 867 -51 925 -17
rect 867 -85 879 -51
rect 913 -85 925 -51
rect 867 -100 925 -85
rect 995 85 1053 100
rect 995 51 1007 85
rect 1041 51 1053 85
rect 995 17 1053 51
rect 995 -17 1007 17
rect 1041 -17 1053 17
rect 995 -51 1053 -17
rect 995 -85 1007 -51
rect 1041 -85 1053 -51
rect 995 -100 1053 -85
rect 1123 85 1181 100
rect 1123 51 1135 85
rect 1169 51 1181 85
rect 1123 17 1181 51
rect 1123 -17 1135 17
rect 1169 -17 1181 17
rect 1123 -51 1181 -17
rect 1123 -85 1135 -51
rect 1169 -85 1181 -51
rect 1123 -100 1181 -85
rect 1251 85 1309 100
rect 1251 51 1263 85
rect 1297 51 1309 85
rect 1251 17 1309 51
rect 1251 -17 1263 17
rect 1297 -17 1309 17
rect 1251 -51 1309 -17
rect 1251 -85 1263 -51
rect 1297 -85 1309 -51
rect 1251 -100 1309 -85
rect 1379 85 1437 100
rect 1379 51 1391 85
rect 1425 51 1437 85
rect 1379 17 1437 51
rect 1379 -17 1391 17
rect 1425 -17 1437 17
rect 1379 -51 1437 -17
rect 1379 -85 1391 -51
rect 1425 -85 1437 -51
rect 1379 -100 1437 -85
rect 1507 85 1565 100
rect 1507 51 1519 85
rect 1553 51 1565 85
rect 1507 17 1565 51
rect 1507 -17 1519 17
rect 1553 -17 1565 17
rect 1507 -51 1565 -17
rect 1507 -85 1519 -51
rect 1553 -85 1565 -51
rect 1507 -100 1565 -85
rect 1635 85 1693 100
rect 1635 51 1647 85
rect 1681 51 1693 85
rect 1635 17 1693 51
rect 1635 -17 1647 17
rect 1681 -17 1693 17
rect 1635 -51 1693 -17
rect 1635 -85 1647 -51
rect 1681 -85 1693 -51
rect 1635 -100 1693 -85
rect 1763 85 1821 100
rect 1763 51 1775 85
rect 1809 51 1821 85
rect 1763 17 1821 51
rect 1763 -17 1775 17
rect 1809 -17 1821 17
rect 1763 -51 1821 -17
rect 1763 -85 1775 -51
rect 1809 -85 1821 -51
rect 1763 -100 1821 -85
rect 1891 85 1949 100
rect 1891 51 1903 85
rect 1937 51 1949 85
rect 1891 17 1949 51
rect 1891 -17 1903 17
rect 1937 -17 1949 17
rect 1891 -51 1949 -17
rect 1891 -85 1903 -51
rect 1937 -85 1949 -51
rect 1891 -100 1949 -85
<< pdiffc >>
rect -1937 51 -1903 85
rect -1937 -17 -1903 17
rect -1937 -85 -1903 -51
rect -1809 51 -1775 85
rect -1809 -17 -1775 17
rect -1809 -85 -1775 -51
rect -1681 51 -1647 85
rect -1681 -17 -1647 17
rect -1681 -85 -1647 -51
rect -1553 51 -1519 85
rect -1553 -17 -1519 17
rect -1553 -85 -1519 -51
rect -1425 51 -1391 85
rect -1425 -17 -1391 17
rect -1425 -85 -1391 -51
rect -1297 51 -1263 85
rect -1297 -17 -1263 17
rect -1297 -85 -1263 -51
rect -1169 51 -1135 85
rect -1169 -17 -1135 17
rect -1169 -85 -1135 -51
rect -1041 51 -1007 85
rect -1041 -17 -1007 17
rect -1041 -85 -1007 -51
rect -913 51 -879 85
rect -913 -17 -879 17
rect -913 -85 -879 -51
rect -785 51 -751 85
rect -785 -17 -751 17
rect -785 -85 -751 -51
rect -657 51 -623 85
rect -657 -17 -623 17
rect -657 -85 -623 -51
rect -529 51 -495 85
rect -529 -17 -495 17
rect -529 -85 -495 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -273 51 -239 85
rect -273 -17 -239 17
rect -273 -85 -239 -51
rect -145 51 -111 85
rect -145 -17 -111 17
rect -145 -85 -111 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 111 51 145 85
rect 111 -17 145 17
rect 111 -85 145 -51
rect 239 51 273 85
rect 239 -17 273 17
rect 239 -85 273 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 495 51 529 85
rect 495 -17 529 17
rect 495 -85 529 -51
rect 623 51 657 85
rect 623 -17 657 17
rect 623 -85 657 -51
rect 751 51 785 85
rect 751 -17 785 17
rect 751 -85 785 -51
rect 879 51 913 85
rect 879 -17 913 17
rect 879 -85 913 -51
rect 1007 51 1041 85
rect 1007 -17 1041 17
rect 1007 -85 1041 -51
rect 1135 51 1169 85
rect 1135 -17 1169 17
rect 1135 -85 1169 -51
rect 1263 51 1297 85
rect 1263 -17 1297 17
rect 1263 -85 1297 -51
rect 1391 51 1425 85
rect 1391 -17 1425 17
rect 1391 -85 1425 -51
rect 1519 51 1553 85
rect 1519 -17 1553 17
rect 1519 -85 1553 -51
rect 1647 51 1681 85
rect 1647 -17 1681 17
rect 1647 -85 1681 -51
rect 1775 51 1809 85
rect 1775 -17 1809 17
rect 1775 -85 1809 -51
rect 1903 51 1937 85
rect 1903 -17 1937 17
rect 1903 -85 1937 -51
<< nsubdiff >>
rect -2051 249 -1955 283
rect -1921 249 -1887 283
rect -1853 249 -1819 283
rect -1785 249 -1751 283
rect -1717 249 -1683 283
rect -1649 249 -1615 283
rect -1581 249 -1547 283
rect -1513 249 -1479 283
rect -1445 249 -1411 283
rect -1377 249 -1343 283
rect -1309 249 -1275 283
rect -1241 249 -1207 283
rect -1173 249 -1139 283
rect -1105 249 -1071 283
rect -1037 249 -1003 283
rect -969 249 -935 283
rect -901 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 901 283
rect 935 249 969 283
rect 1003 249 1037 283
rect 1071 249 1105 283
rect 1139 249 1173 283
rect 1207 249 1241 283
rect 1275 249 1309 283
rect 1343 249 1377 283
rect 1411 249 1445 283
rect 1479 249 1513 283
rect 1547 249 1581 283
rect 1615 249 1649 283
rect 1683 249 1717 283
rect 1751 249 1785 283
rect 1819 249 1853 283
rect 1887 249 1921 283
rect 1955 249 2051 283
rect -2051 187 -2017 249
rect -2051 119 -2017 153
rect 2017 187 2051 249
rect 2017 119 2051 153
rect -2051 51 -2017 85
rect -2051 -17 -2017 17
rect -2051 -85 -2017 -51
rect 2017 51 2051 85
rect 2017 -17 2051 17
rect 2017 -85 2051 -51
rect -2051 -153 -2017 -119
rect -2051 -249 -2017 -187
rect 2017 -153 2051 -119
rect 2017 -249 2051 -187
rect -2051 -283 -1955 -249
rect -1921 -283 -1887 -249
rect -1853 -283 -1819 -249
rect -1785 -283 -1751 -249
rect -1717 -283 -1683 -249
rect -1649 -283 -1615 -249
rect -1581 -283 -1547 -249
rect -1513 -283 -1479 -249
rect -1445 -283 -1411 -249
rect -1377 -283 -1343 -249
rect -1309 -283 -1275 -249
rect -1241 -283 -1207 -249
rect -1173 -283 -1139 -249
rect -1105 -283 -1071 -249
rect -1037 -283 -1003 -249
rect -969 -283 -935 -249
rect -901 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 901 -249
rect 935 -283 969 -249
rect 1003 -283 1037 -249
rect 1071 -283 1105 -249
rect 1139 -283 1173 -249
rect 1207 -283 1241 -249
rect 1275 -283 1309 -249
rect 1343 -283 1377 -249
rect 1411 -283 1445 -249
rect 1479 -283 1513 -249
rect 1547 -283 1581 -249
rect 1615 -283 1649 -249
rect 1683 -283 1717 -249
rect 1751 -283 1785 -249
rect 1819 -283 1853 -249
rect 1887 -283 1921 -249
rect 1955 -283 2051 -249
<< nsubdiffcont >>
rect -1955 249 -1921 283
rect -1887 249 -1853 283
rect -1819 249 -1785 283
rect -1751 249 -1717 283
rect -1683 249 -1649 283
rect -1615 249 -1581 283
rect -1547 249 -1513 283
rect -1479 249 -1445 283
rect -1411 249 -1377 283
rect -1343 249 -1309 283
rect -1275 249 -1241 283
rect -1207 249 -1173 283
rect -1139 249 -1105 283
rect -1071 249 -1037 283
rect -1003 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1003 283
rect 1037 249 1071 283
rect 1105 249 1139 283
rect 1173 249 1207 283
rect 1241 249 1275 283
rect 1309 249 1343 283
rect 1377 249 1411 283
rect 1445 249 1479 283
rect 1513 249 1547 283
rect 1581 249 1615 283
rect 1649 249 1683 283
rect 1717 249 1751 283
rect 1785 249 1819 283
rect 1853 249 1887 283
rect 1921 249 1955 283
rect -2051 153 -2017 187
rect -2051 85 -2017 119
rect 2017 153 2051 187
rect -2051 17 -2017 51
rect -2051 -51 -2017 -17
rect -2051 -119 -2017 -85
rect 2017 85 2051 119
rect 2017 17 2051 51
rect 2017 -51 2051 -17
rect -2051 -187 -2017 -153
rect 2017 -119 2051 -85
rect 2017 -187 2051 -153
rect -1955 -283 -1921 -249
rect -1887 -283 -1853 -249
rect -1819 -283 -1785 -249
rect -1751 -283 -1717 -249
rect -1683 -283 -1649 -249
rect -1615 -283 -1581 -249
rect -1547 -283 -1513 -249
rect -1479 -283 -1445 -249
rect -1411 -283 -1377 -249
rect -1343 -283 -1309 -249
rect -1275 -283 -1241 -249
rect -1207 -283 -1173 -249
rect -1139 -283 -1105 -249
rect -1071 -283 -1037 -249
rect -1003 -283 -969 -249
rect -935 -283 -901 -249
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
rect 901 -283 935 -249
rect 969 -283 1003 -249
rect 1037 -283 1071 -249
rect 1105 -283 1139 -249
rect 1173 -283 1207 -249
rect 1241 -283 1275 -249
rect 1309 -283 1343 -249
rect 1377 -283 1411 -249
rect 1445 -283 1479 -249
rect 1513 -283 1547 -249
rect 1581 -283 1615 -249
rect 1649 -283 1683 -249
rect 1717 -283 1751 -249
rect 1785 -283 1819 -249
rect 1853 -283 1887 -249
rect 1921 -283 1955 -249
<< poly >>
rect -1891 181 -1821 197
rect -1891 147 -1873 181
rect -1839 147 -1821 181
rect -1891 100 -1821 147
rect -1763 181 -1693 197
rect -1763 147 -1745 181
rect -1711 147 -1693 181
rect -1763 100 -1693 147
rect -1635 181 -1565 197
rect -1635 147 -1617 181
rect -1583 147 -1565 181
rect -1635 100 -1565 147
rect -1507 181 -1437 197
rect -1507 147 -1489 181
rect -1455 147 -1437 181
rect -1507 100 -1437 147
rect -1379 181 -1309 197
rect -1379 147 -1361 181
rect -1327 147 -1309 181
rect -1379 100 -1309 147
rect -1251 181 -1181 197
rect -1251 147 -1233 181
rect -1199 147 -1181 181
rect -1251 100 -1181 147
rect -1123 181 -1053 197
rect -1123 147 -1105 181
rect -1071 147 -1053 181
rect -1123 100 -1053 147
rect -995 181 -925 197
rect -995 147 -977 181
rect -943 147 -925 181
rect -995 100 -925 147
rect -867 181 -797 197
rect -867 147 -849 181
rect -815 147 -797 181
rect -867 100 -797 147
rect -739 181 -669 197
rect -739 147 -721 181
rect -687 147 -669 181
rect -739 100 -669 147
rect -611 181 -541 197
rect -611 147 -593 181
rect -559 147 -541 181
rect -611 100 -541 147
rect -483 181 -413 197
rect -483 147 -465 181
rect -431 147 -413 181
rect -483 100 -413 147
rect -355 181 -285 197
rect -355 147 -337 181
rect -303 147 -285 181
rect -355 100 -285 147
rect -227 181 -157 197
rect -227 147 -209 181
rect -175 147 -157 181
rect -227 100 -157 147
rect -99 181 -29 197
rect -99 147 -81 181
rect -47 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 47 181
rect 81 147 99 181
rect 29 100 99 147
rect 157 181 227 197
rect 157 147 175 181
rect 209 147 227 181
rect 157 100 227 147
rect 285 181 355 197
rect 285 147 303 181
rect 337 147 355 181
rect 285 100 355 147
rect 413 181 483 197
rect 413 147 431 181
rect 465 147 483 181
rect 413 100 483 147
rect 541 181 611 197
rect 541 147 559 181
rect 593 147 611 181
rect 541 100 611 147
rect 669 181 739 197
rect 669 147 687 181
rect 721 147 739 181
rect 669 100 739 147
rect 797 181 867 197
rect 797 147 815 181
rect 849 147 867 181
rect 797 100 867 147
rect 925 181 995 197
rect 925 147 943 181
rect 977 147 995 181
rect 925 100 995 147
rect 1053 181 1123 197
rect 1053 147 1071 181
rect 1105 147 1123 181
rect 1053 100 1123 147
rect 1181 181 1251 197
rect 1181 147 1199 181
rect 1233 147 1251 181
rect 1181 100 1251 147
rect 1309 181 1379 197
rect 1309 147 1327 181
rect 1361 147 1379 181
rect 1309 100 1379 147
rect 1437 181 1507 197
rect 1437 147 1455 181
rect 1489 147 1507 181
rect 1437 100 1507 147
rect 1565 181 1635 197
rect 1565 147 1583 181
rect 1617 147 1635 181
rect 1565 100 1635 147
rect 1693 181 1763 197
rect 1693 147 1711 181
rect 1745 147 1763 181
rect 1693 100 1763 147
rect 1821 181 1891 197
rect 1821 147 1839 181
rect 1873 147 1891 181
rect 1821 100 1891 147
rect -1891 -147 -1821 -100
rect -1891 -181 -1873 -147
rect -1839 -181 -1821 -147
rect -1891 -197 -1821 -181
rect -1763 -147 -1693 -100
rect -1763 -181 -1745 -147
rect -1711 -181 -1693 -147
rect -1763 -197 -1693 -181
rect -1635 -147 -1565 -100
rect -1635 -181 -1617 -147
rect -1583 -181 -1565 -147
rect -1635 -197 -1565 -181
rect -1507 -147 -1437 -100
rect -1507 -181 -1489 -147
rect -1455 -181 -1437 -147
rect -1507 -197 -1437 -181
rect -1379 -147 -1309 -100
rect -1379 -181 -1361 -147
rect -1327 -181 -1309 -147
rect -1379 -197 -1309 -181
rect -1251 -147 -1181 -100
rect -1251 -181 -1233 -147
rect -1199 -181 -1181 -147
rect -1251 -197 -1181 -181
rect -1123 -147 -1053 -100
rect -1123 -181 -1105 -147
rect -1071 -181 -1053 -147
rect -1123 -197 -1053 -181
rect -995 -147 -925 -100
rect -995 -181 -977 -147
rect -943 -181 -925 -147
rect -995 -197 -925 -181
rect -867 -147 -797 -100
rect -867 -181 -849 -147
rect -815 -181 -797 -147
rect -867 -197 -797 -181
rect -739 -147 -669 -100
rect -739 -181 -721 -147
rect -687 -181 -669 -147
rect -739 -197 -669 -181
rect -611 -147 -541 -100
rect -611 -181 -593 -147
rect -559 -181 -541 -147
rect -611 -197 -541 -181
rect -483 -147 -413 -100
rect -483 -181 -465 -147
rect -431 -181 -413 -147
rect -483 -197 -413 -181
rect -355 -147 -285 -100
rect -355 -181 -337 -147
rect -303 -181 -285 -147
rect -355 -197 -285 -181
rect -227 -147 -157 -100
rect -227 -181 -209 -147
rect -175 -181 -157 -147
rect -227 -197 -157 -181
rect -99 -147 -29 -100
rect -99 -181 -81 -147
rect -47 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 47 -147
rect 81 -181 99 -147
rect 29 -197 99 -181
rect 157 -147 227 -100
rect 157 -181 175 -147
rect 209 -181 227 -147
rect 157 -197 227 -181
rect 285 -147 355 -100
rect 285 -181 303 -147
rect 337 -181 355 -147
rect 285 -197 355 -181
rect 413 -147 483 -100
rect 413 -181 431 -147
rect 465 -181 483 -147
rect 413 -197 483 -181
rect 541 -147 611 -100
rect 541 -181 559 -147
rect 593 -181 611 -147
rect 541 -197 611 -181
rect 669 -147 739 -100
rect 669 -181 687 -147
rect 721 -181 739 -147
rect 669 -197 739 -181
rect 797 -147 867 -100
rect 797 -181 815 -147
rect 849 -181 867 -147
rect 797 -197 867 -181
rect 925 -147 995 -100
rect 925 -181 943 -147
rect 977 -181 995 -147
rect 925 -197 995 -181
rect 1053 -147 1123 -100
rect 1053 -181 1071 -147
rect 1105 -181 1123 -147
rect 1053 -197 1123 -181
rect 1181 -147 1251 -100
rect 1181 -181 1199 -147
rect 1233 -181 1251 -147
rect 1181 -197 1251 -181
rect 1309 -147 1379 -100
rect 1309 -181 1327 -147
rect 1361 -181 1379 -147
rect 1309 -197 1379 -181
rect 1437 -147 1507 -100
rect 1437 -181 1455 -147
rect 1489 -181 1507 -147
rect 1437 -197 1507 -181
rect 1565 -147 1635 -100
rect 1565 -181 1583 -147
rect 1617 -181 1635 -147
rect 1565 -197 1635 -181
rect 1693 -147 1763 -100
rect 1693 -181 1711 -147
rect 1745 -181 1763 -147
rect 1693 -197 1763 -181
rect 1821 -147 1891 -100
rect 1821 -181 1839 -147
rect 1873 -181 1891 -147
rect 1821 -197 1891 -181
<< polycont >>
rect -1873 147 -1839 181
rect -1745 147 -1711 181
rect -1617 147 -1583 181
rect -1489 147 -1455 181
rect -1361 147 -1327 181
rect -1233 147 -1199 181
rect -1105 147 -1071 181
rect -977 147 -943 181
rect -849 147 -815 181
rect -721 147 -687 181
rect -593 147 -559 181
rect -465 147 -431 181
rect -337 147 -303 181
rect -209 147 -175 181
rect -81 147 -47 181
rect 47 147 81 181
rect 175 147 209 181
rect 303 147 337 181
rect 431 147 465 181
rect 559 147 593 181
rect 687 147 721 181
rect 815 147 849 181
rect 943 147 977 181
rect 1071 147 1105 181
rect 1199 147 1233 181
rect 1327 147 1361 181
rect 1455 147 1489 181
rect 1583 147 1617 181
rect 1711 147 1745 181
rect 1839 147 1873 181
rect -1873 -181 -1839 -147
rect -1745 -181 -1711 -147
rect -1617 -181 -1583 -147
rect -1489 -181 -1455 -147
rect -1361 -181 -1327 -147
rect -1233 -181 -1199 -147
rect -1105 -181 -1071 -147
rect -977 -181 -943 -147
rect -849 -181 -815 -147
rect -721 -181 -687 -147
rect -593 -181 -559 -147
rect -465 -181 -431 -147
rect -337 -181 -303 -147
rect -209 -181 -175 -147
rect -81 -181 -47 -147
rect 47 -181 81 -147
rect 175 -181 209 -147
rect 303 -181 337 -147
rect 431 -181 465 -147
rect 559 -181 593 -147
rect 687 -181 721 -147
rect 815 -181 849 -147
rect 943 -181 977 -147
rect 1071 -181 1105 -147
rect 1199 -181 1233 -147
rect 1327 -181 1361 -147
rect 1455 -181 1489 -147
rect 1583 -181 1617 -147
rect 1711 -181 1745 -147
rect 1839 -181 1873 -147
<< locali >>
rect -2051 249 -1955 283
rect -1921 249 -1887 283
rect -1853 249 -1819 283
rect -1785 249 -1751 283
rect -1717 249 -1683 283
rect -1649 249 -1615 283
rect -1581 249 -1547 283
rect -1513 249 -1479 283
rect -1445 249 -1411 283
rect -1377 249 -1343 283
rect -1309 249 -1275 283
rect -1241 249 -1207 283
rect -1173 249 -1139 283
rect -1105 249 -1071 283
rect -1037 249 -1003 283
rect -969 249 -935 283
rect -901 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 901 283
rect 935 249 969 283
rect 1003 249 1037 283
rect 1071 249 1105 283
rect 1139 249 1173 283
rect 1207 249 1241 283
rect 1275 249 1309 283
rect 1343 249 1377 283
rect 1411 249 1445 283
rect 1479 249 1513 283
rect 1547 249 1581 283
rect 1615 249 1649 283
rect 1683 249 1717 283
rect 1751 249 1785 283
rect 1819 249 1853 283
rect 1887 249 1921 283
rect 1955 249 2051 283
rect -2051 187 -2017 249
rect 2017 187 2051 249
rect -2051 119 -2017 153
rect -1891 147 -1873 181
rect -1839 147 -1821 181
rect -1763 147 -1745 181
rect -1711 147 -1693 181
rect -1635 147 -1617 181
rect -1583 147 -1565 181
rect -1507 147 -1489 181
rect -1455 147 -1437 181
rect -1379 147 -1361 181
rect -1327 147 -1309 181
rect -1251 147 -1233 181
rect -1199 147 -1181 181
rect -1123 147 -1105 181
rect -1071 147 -1053 181
rect -995 147 -977 181
rect -943 147 -925 181
rect -867 147 -849 181
rect -815 147 -797 181
rect -739 147 -721 181
rect -687 147 -669 181
rect -611 147 -593 181
rect -559 147 -541 181
rect -483 147 -465 181
rect -431 147 -413 181
rect -355 147 -337 181
rect -303 147 -285 181
rect -227 147 -209 181
rect -175 147 -157 181
rect -99 147 -81 181
rect -47 147 -29 181
rect 29 147 47 181
rect 81 147 99 181
rect 157 147 175 181
rect 209 147 227 181
rect 285 147 303 181
rect 337 147 355 181
rect 413 147 431 181
rect 465 147 483 181
rect 541 147 559 181
rect 593 147 611 181
rect 669 147 687 181
rect 721 147 739 181
rect 797 147 815 181
rect 849 147 867 181
rect 925 147 943 181
rect 977 147 995 181
rect 1053 147 1071 181
rect 1105 147 1123 181
rect 1181 147 1199 181
rect 1233 147 1251 181
rect 1309 147 1327 181
rect 1361 147 1379 181
rect 1437 147 1455 181
rect 1489 147 1507 181
rect 1565 147 1583 181
rect 1617 147 1635 181
rect 1693 147 1711 181
rect 1745 147 1763 181
rect 1821 147 1839 181
rect 1873 147 1891 181
rect 2017 119 2051 153
rect -2051 51 -2017 85
rect -2051 -17 -2017 17
rect -2051 -85 -2017 -51
rect -1937 85 -1903 104
rect -1937 17 -1903 19
rect -1937 -19 -1903 -17
rect -1937 -104 -1903 -85
rect -1809 85 -1775 104
rect -1809 17 -1775 19
rect -1809 -19 -1775 -17
rect -1809 -104 -1775 -85
rect -1681 85 -1647 104
rect -1681 17 -1647 19
rect -1681 -19 -1647 -17
rect -1681 -104 -1647 -85
rect -1553 85 -1519 104
rect -1553 17 -1519 19
rect -1553 -19 -1519 -17
rect -1553 -104 -1519 -85
rect -1425 85 -1391 104
rect -1425 17 -1391 19
rect -1425 -19 -1391 -17
rect -1425 -104 -1391 -85
rect -1297 85 -1263 104
rect -1297 17 -1263 19
rect -1297 -19 -1263 -17
rect -1297 -104 -1263 -85
rect -1169 85 -1135 104
rect -1169 17 -1135 19
rect -1169 -19 -1135 -17
rect -1169 -104 -1135 -85
rect -1041 85 -1007 104
rect -1041 17 -1007 19
rect -1041 -19 -1007 -17
rect -1041 -104 -1007 -85
rect -913 85 -879 104
rect -913 17 -879 19
rect -913 -19 -879 -17
rect -913 -104 -879 -85
rect -785 85 -751 104
rect -785 17 -751 19
rect -785 -19 -751 -17
rect -785 -104 -751 -85
rect -657 85 -623 104
rect -657 17 -623 19
rect -657 -19 -623 -17
rect -657 -104 -623 -85
rect -529 85 -495 104
rect -529 17 -495 19
rect -529 -19 -495 -17
rect -529 -104 -495 -85
rect -401 85 -367 104
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -104 -367 -85
rect -273 85 -239 104
rect -273 17 -239 19
rect -273 -19 -239 -17
rect -273 -104 -239 -85
rect -145 85 -111 104
rect -145 17 -111 19
rect -145 -19 -111 -17
rect -145 -104 -111 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 111 85 145 104
rect 111 17 145 19
rect 111 -19 145 -17
rect 111 -104 145 -85
rect 239 85 273 104
rect 239 17 273 19
rect 239 -19 273 -17
rect 239 -104 273 -85
rect 367 85 401 104
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -104 401 -85
rect 495 85 529 104
rect 495 17 529 19
rect 495 -19 529 -17
rect 495 -104 529 -85
rect 623 85 657 104
rect 623 17 657 19
rect 623 -19 657 -17
rect 623 -104 657 -85
rect 751 85 785 104
rect 751 17 785 19
rect 751 -19 785 -17
rect 751 -104 785 -85
rect 879 85 913 104
rect 879 17 913 19
rect 879 -19 913 -17
rect 879 -104 913 -85
rect 1007 85 1041 104
rect 1007 17 1041 19
rect 1007 -19 1041 -17
rect 1007 -104 1041 -85
rect 1135 85 1169 104
rect 1135 17 1169 19
rect 1135 -19 1169 -17
rect 1135 -104 1169 -85
rect 1263 85 1297 104
rect 1263 17 1297 19
rect 1263 -19 1297 -17
rect 1263 -104 1297 -85
rect 1391 85 1425 104
rect 1391 17 1425 19
rect 1391 -19 1425 -17
rect 1391 -104 1425 -85
rect 1519 85 1553 104
rect 1519 17 1553 19
rect 1519 -19 1553 -17
rect 1519 -104 1553 -85
rect 1647 85 1681 104
rect 1647 17 1681 19
rect 1647 -19 1681 -17
rect 1647 -104 1681 -85
rect 1775 85 1809 104
rect 1775 17 1809 19
rect 1775 -19 1809 -17
rect 1775 -104 1809 -85
rect 1903 85 1937 104
rect 1903 17 1937 19
rect 1903 -19 1937 -17
rect 1903 -104 1937 -85
rect 2017 51 2051 85
rect 2017 -17 2051 17
rect 2017 -85 2051 -51
rect -2051 -153 -2017 -119
rect -1891 -181 -1873 -147
rect -1839 -181 -1821 -147
rect -1763 -181 -1745 -147
rect -1711 -181 -1693 -147
rect -1635 -181 -1617 -147
rect -1583 -181 -1565 -147
rect -1507 -181 -1489 -147
rect -1455 -181 -1437 -147
rect -1379 -181 -1361 -147
rect -1327 -181 -1309 -147
rect -1251 -181 -1233 -147
rect -1199 -181 -1181 -147
rect -1123 -181 -1105 -147
rect -1071 -181 -1053 -147
rect -995 -181 -977 -147
rect -943 -181 -925 -147
rect -867 -181 -849 -147
rect -815 -181 -797 -147
rect -739 -181 -721 -147
rect -687 -181 -669 -147
rect -611 -181 -593 -147
rect -559 -181 -541 -147
rect -483 -181 -465 -147
rect -431 -181 -413 -147
rect -355 -181 -337 -147
rect -303 -181 -285 -147
rect -227 -181 -209 -147
rect -175 -181 -157 -147
rect -99 -181 -81 -147
rect -47 -181 -29 -147
rect 29 -181 47 -147
rect 81 -181 99 -147
rect 157 -181 175 -147
rect 209 -181 227 -147
rect 285 -181 303 -147
rect 337 -181 355 -147
rect 413 -181 431 -147
rect 465 -181 483 -147
rect 541 -181 559 -147
rect 593 -181 611 -147
rect 669 -181 687 -147
rect 721 -181 739 -147
rect 797 -181 815 -147
rect 849 -181 867 -147
rect 925 -181 943 -147
rect 977 -181 995 -147
rect 1053 -181 1071 -147
rect 1105 -181 1123 -147
rect 1181 -181 1199 -147
rect 1233 -181 1251 -147
rect 1309 -181 1327 -147
rect 1361 -181 1379 -147
rect 1437 -181 1455 -147
rect 1489 -181 1507 -147
rect 1565 -181 1583 -147
rect 1617 -181 1635 -147
rect 1693 -181 1711 -147
rect 1745 -181 1763 -147
rect 1821 -181 1839 -147
rect 1873 -181 1891 -147
rect 2017 -153 2051 -119
rect -2051 -249 -2017 -187
rect 2017 -249 2051 -187
rect -2051 -283 -1955 -249
rect -1921 -283 -1887 -249
rect -1853 -283 -1819 -249
rect -1785 -283 -1751 -249
rect -1717 -283 -1683 -249
rect -1649 -283 -1615 -249
rect -1581 -283 -1547 -249
rect -1513 -283 -1479 -249
rect -1445 -283 -1411 -249
rect -1377 -283 -1343 -249
rect -1309 -283 -1275 -249
rect -1241 -283 -1207 -249
rect -1173 -283 -1139 -249
rect -1105 -283 -1071 -249
rect -1037 -283 -1003 -249
rect -969 -283 -935 -249
rect -901 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 901 -249
rect 935 -283 969 -249
rect 1003 -283 1037 -249
rect 1071 -283 1105 -249
rect 1139 -283 1173 -249
rect 1207 -283 1241 -249
rect 1275 -283 1309 -249
rect 1343 -283 1377 -249
rect 1411 -283 1445 -249
rect 1479 -283 1513 -249
rect 1547 -283 1581 -249
rect 1615 -283 1649 -249
rect 1683 -283 1717 -249
rect 1751 -283 1785 -249
rect 1819 -283 1853 -249
rect 1887 -283 1921 -249
rect 1955 -283 2051 -249
<< viali >>
rect -1873 147 -1839 181
rect -1745 147 -1711 181
rect -1617 147 -1583 181
rect -1489 147 -1455 181
rect -1361 147 -1327 181
rect -1233 147 -1199 181
rect -1105 147 -1071 181
rect -977 147 -943 181
rect -849 147 -815 181
rect -721 147 -687 181
rect -593 147 -559 181
rect -465 147 -431 181
rect -337 147 -303 181
rect -209 147 -175 181
rect -81 147 -47 181
rect 47 147 81 181
rect 175 147 209 181
rect 303 147 337 181
rect 431 147 465 181
rect 559 147 593 181
rect 687 147 721 181
rect 815 147 849 181
rect 943 147 977 181
rect 1071 147 1105 181
rect 1199 147 1233 181
rect 1327 147 1361 181
rect 1455 147 1489 181
rect 1583 147 1617 181
rect 1711 147 1745 181
rect 1839 147 1873 181
rect -1937 51 -1903 53
rect -1937 19 -1903 51
rect -1937 -51 -1903 -19
rect -1937 -53 -1903 -51
rect -1809 51 -1775 53
rect -1809 19 -1775 51
rect -1809 -51 -1775 -19
rect -1809 -53 -1775 -51
rect -1681 51 -1647 53
rect -1681 19 -1647 51
rect -1681 -51 -1647 -19
rect -1681 -53 -1647 -51
rect -1553 51 -1519 53
rect -1553 19 -1519 51
rect -1553 -51 -1519 -19
rect -1553 -53 -1519 -51
rect -1425 51 -1391 53
rect -1425 19 -1391 51
rect -1425 -51 -1391 -19
rect -1425 -53 -1391 -51
rect -1297 51 -1263 53
rect -1297 19 -1263 51
rect -1297 -51 -1263 -19
rect -1297 -53 -1263 -51
rect -1169 51 -1135 53
rect -1169 19 -1135 51
rect -1169 -51 -1135 -19
rect -1169 -53 -1135 -51
rect -1041 51 -1007 53
rect -1041 19 -1007 51
rect -1041 -51 -1007 -19
rect -1041 -53 -1007 -51
rect -913 51 -879 53
rect -913 19 -879 51
rect -913 -51 -879 -19
rect -913 -53 -879 -51
rect -785 51 -751 53
rect -785 19 -751 51
rect -785 -51 -751 -19
rect -785 -53 -751 -51
rect -657 51 -623 53
rect -657 19 -623 51
rect -657 -51 -623 -19
rect -657 -53 -623 -51
rect -529 51 -495 53
rect -529 19 -495 51
rect -529 -51 -495 -19
rect -529 -53 -495 -51
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -273 51 -239 53
rect -273 19 -239 51
rect -273 -51 -239 -19
rect -273 -53 -239 -51
rect -145 51 -111 53
rect -145 19 -111 51
rect -145 -51 -111 -19
rect -145 -53 -111 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 111 51 145 53
rect 111 19 145 51
rect 111 -51 145 -19
rect 111 -53 145 -51
rect 239 51 273 53
rect 239 19 273 51
rect 239 -51 273 -19
rect 239 -53 273 -51
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 495 51 529 53
rect 495 19 529 51
rect 495 -51 529 -19
rect 495 -53 529 -51
rect 623 51 657 53
rect 623 19 657 51
rect 623 -51 657 -19
rect 623 -53 657 -51
rect 751 51 785 53
rect 751 19 785 51
rect 751 -51 785 -19
rect 751 -53 785 -51
rect 879 51 913 53
rect 879 19 913 51
rect 879 -51 913 -19
rect 879 -53 913 -51
rect 1007 51 1041 53
rect 1007 19 1041 51
rect 1007 -51 1041 -19
rect 1007 -53 1041 -51
rect 1135 51 1169 53
rect 1135 19 1169 51
rect 1135 -51 1169 -19
rect 1135 -53 1169 -51
rect 1263 51 1297 53
rect 1263 19 1297 51
rect 1263 -51 1297 -19
rect 1263 -53 1297 -51
rect 1391 51 1425 53
rect 1391 19 1425 51
rect 1391 -51 1425 -19
rect 1391 -53 1425 -51
rect 1519 51 1553 53
rect 1519 19 1553 51
rect 1519 -51 1553 -19
rect 1519 -53 1553 -51
rect 1647 51 1681 53
rect 1647 19 1681 51
rect 1647 -51 1681 -19
rect 1647 -53 1681 -51
rect 1775 51 1809 53
rect 1775 19 1809 51
rect 1775 -51 1809 -19
rect 1775 -53 1809 -51
rect 1903 51 1937 53
rect 1903 19 1937 51
rect 1903 -51 1937 -19
rect 1903 -53 1937 -51
rect -1873 -181 -1839 -147
rect -1745 -181 -1711 -147
rect -1617 -181 -1583 -147
rect -1489 -181 -1455 -147
rect -1361 -181 -1327 -147
rect -1233 -181 -1199 -147
rect -1105 -181 -1071 -147
rect -977 -181 -943 -147
rect -849 -181 -815 -147
rect -721 -181 -687 -147
rect -593 -181 -559 -147
rect -465 -181 -431 -147
rect -337 -181 -303 -147
rect -209 -181 -175 -147
rect -81 -181 -47 -147
rect 47 -181 81 -147
rect 175 -181 209 -147
rect 303 -181 337 -147
rect 431 -181 465 -147
rect 559 -181 593 -147
rect 687 -181 721 -147
rect 815 -181 849 -147
rect 943 -181 977 -147
rect 1071 -181 1105 -147
rect 1199 -181 1233 -147
rect 1327 -181 1361 -147
rect 1455 -181 1489 -147
rect 1583 -181 1617 -147
rect 1711 -181 1745 -147
rect 1839 -181 1873 -147
<< metal1 >>
rect -1887 181 -1825 187
rect -1887 147 -1873 181
rect -1839 147 -1825 181
rect -1887 141 -1825 147
rect -1759 181 -1697 187
rect -1759 147 -1745 181
rect -1711 147 -1697 181
rect -1759 141 -1697 147
rect -1631 181 -1569 187
rect -1631 147 -1617 181
rect -1583 147 -1569 181
rect -1631 141 -1569 147
rect -1503 181 -1441 187
rect -1503 147 -1489 181
rect -1455 147 -1441 181
rect -1503 141 -1441 147
rect -1375 181 -1313 187
rect -1375 147 -1361 181
rect -1327 147 -1313 181
rect -1375 141 -1313 147
rect -1247 181 -1185 187
rect -1247 147 -1233 181
rect -1199 147 -1185 181
rect -1247 141 -1185 147
rect -1119 181 -1057 187
rect -1119 147 -1105 181
rect -1071 147 -1057 181
rect -1119 141 -1057 147
rect -991 181 -929 187
rect -991 147 -977 181
rect -943 147 -929 181
rect -991 141 -929 147
rect -863 181 -801 187
rect -863 147 -849 181
rect -815 147 -801 181
rect -863 141 -801 147
rect -735 181 -673 187
rect -735 147 -721 181
rect -687 147 -673 181
rect -735 141 -673 147
rect -607 181 -545 187
rect -607 147 -593 181
rect -559 147 -545 181
rect -607 141 -545 147
rect -479 181 -417 187
rect -479 147 -465 181
rect -431 147 -417 181
rect -479 141 -417 147
rect -351 181 -289 187
rect -351 147 -337 181
rect -303 147 -289 181
rect -351 141 -289 147
rect -223 181 -161 187
rect -223 147 -209 181
rect -175 147 -161 181
rect -223 141 -161 147
rect -95 181 -33 187
rect -95 147 -81 181
rect -47 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 47 181
rect 81 147 95 181
rect 33 141 95 147
rect 161 181 223 187
rect 161 147 175 181
rect 209 147 223 181
rect 161 141 223 147
rect 289 181 351 187
rect 289 147 303 181
rect 337 147 351 181
rect 289 141 351 147
rect 417 181 479 187
rect 417 147 431 181
rect 465 147 479 181
rect 417 141 479 147
rect 545 181 607 187
rect 545 147 559 181
rect 593 147 607 181
rect 545 141 607 147
rect 673 181 735 187
rect 673 147 687 181
rect 721 147 735 181
rect 673 141 735 147
rect 801 181 863 187
rect 801 147 815 181
rect 849 147 863 181
rect 801 141 863 147
rect 929 181 991 187
rect 929 147 943 181
rect 977 147 991 181
rect 929 141 991 147
rect 1057 181 1119 187
rect 1057 147 1071 181
rect 1105 147 1119 181
rect 1057 141 1119 147
rect 1185 181 1247 187
rect 1185 147 1199 181
rect 1233 147 1247 181
rect 1185 141 1247 147
rect 1313 181 1375 187
rect 1313 147 1327 181
rect 1361 147 1375 181
rect 1313 141 1375 147
rect 1441 181 1503 187
rect 1441 147 1455 181
rect 1489 147 1503 181
rect 1441 141 1503 147
rect 1569 181 1631 187
rect 1569 147 1583 181
rect 1617 147 1631 181
rect 1569 141 1631 147
rect 1697 181 1759 187
rect 1697 147 1711 181
rect 1745 147 1759 181
rect 1697 141 1759 147
rect 1825 181 1887 187
rect 1825 147 1839 181
rect 1873 147 1887 181
rect 1825 141 1887 147
rect -1943 53 -1897 100
rect -1943 19 -1937 53
rect -1903 19 -1897 53
rect -1943 -19 -1897 19
rect -1943 -53 -1937 -19
rect -1903 -53 -1897 -19
rect -1943 -100 -1897 -53
rect -1815 53 -1769 100
rect -1815 19 -1809 53
rect -1775 19 -1769 53
rect -1815 -19 -1769 19
rect -1815 -53 -1809 -19
rect -1775 -53 -1769 -19
rect -1815 -100 -1769 -53
rect -1687 53 -1641 100
rect -1687 19 -1681 53
rect -1647 19 -1641 53
rect -1687 -19 -1641 19
rect -1687 -53 -1681 -19
rect -1647 -53 -1641 -19
rect -1687 -100 -1641 -53
rect -1559 53 -1513 100
rect -1559 19 -1553 53
rect -1519 19 -1513 53
rect -1559 -19 -1513 19
rect -1559 -53 -1553 -19
rect -1519 -53 -1513 -19
rect -1559 -100 -1513 -53
rect -1431 53 -1385 100
rect -1431 19 -1425 53
rect -1391 19 -1385 53
rect -1431 -19 -1385 19
rect -1431 -53 -1425 -19
rect -1391 -53 -1385 -19
rect -1431 -100 -1385 -53
rect -1303 53 -1257 100
rect -1303 19 -1297 53
rect -1263 19 -1257 53
rect -1303 -19 -1257 19
rect -1303 -53 -1297 -19
rect -1263 -53 -1257 -19
rect -1303 -100 -1257 -53
rect -1175 53 -1129 100
rect -1175 19 -1169 53
rect -1135 19 -1129 53
rect -1175 -19 -1129 19
rect -1175 -53 -1169 -19
rect -1135 -53 -1129 -19
rect -1175 -100 -1129 -53
rect -1047 53 -1001 100
rect -1047 19 -1041 53
rect -1007 19 -1001 53
rect -1047 -19 -1001 19
rect -1047 -53 -1041 -19
rect -1007 -53 -1001 -19
rect -1047 -100 -1001 -53
rect -919 53 -873 100
rect -919 19 -913 53
rect -879 19 -873 53
rect -919 -19 -873 19
rect -919 -53 -913 -19
rect -879 -53 -873 -19
rect -919 -100 -873 -53
rect -791 53 -745 100
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -100 -745 -53
rect -663 53 -617 100
rect -663 19 -657 53
rect -623 19 -617 53
rect -663 -19 -617 19
rect -663 -53 -657 -19
rect -623 -53 -617 -19
rect -663 -100 -617 -53
rect -535 53 -489 100
rect -535 19 -529 53
rect -495 19 -489 53
rect -535 -19 -489 19
rect -535 -53 -529 -19
rect -495 -53 -489 -19
rect -535 -100 -489 -53
rect -407 53 -361 100
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -100 -361 -53
rect -279 53 -233 100
rect -279 19 -273 53
rect -239 19 -233 53
rect -279 -19 -233 19
rect -279 -53 -273 -19
rect -239 -53 -233 -19
rect -279 -100 -233 -53
rect -151 53 -105 100
rect -151 19 -145 53
rect -111 19 -105 53
rect -151 -19 -105 19
rect -151 -53 -145 -19
rect -111 -53 -105 -19
rect -151 -100 -105 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 105 53 151 100
rect 105 19 111 53
rect 145 19 151 53
rect 105 -19 151 19
rect 105 -53 111 -19
rect 145 -53 151 -19
rect 105 -100 151 -53
rect 233 53 279 100
rect 233 19 239 53
rect 273 19 279 53
rect 233 -19 279 19
rect 233 -53 239 -19
rect 273 -53 279 -19
rect 233 -100 279 -53
rect 361 53 407 100
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -100 407 -53
rect 489 53 535 100
rect 489 19 495 53
rect 529 19 535 53
rect 489 -19 535 19
rect 489 -53 495 -19
rect 529 -53 535 -19
rect 489 -100 535 -53
rect 617 53 663 100
rect 617 19 623 53
rect 657 19 663 53
rect 617 -19 663 19
rect 617 -53 623 -19
rect 657 -53 663 -19
rect 617 -100 663 -53
rect 745 53 791 100
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -100 791 -53
rect 873 53 919 100
rect 873 19 879 53
rect 913 19 919 53
rect 873 -19 919 19
rect 873 -53 879 -19
rect 913 -53 919 -19
rect 873 -100 919 -53
rect 1001 53 1047 100
rect 1001 19 1007 53
rect 1041 19 1047 53
rect 1001 -19 1047 19
rect 1001 -53 1007 -19
rect 1041 -53 1047 -19
rect 1001 -100 1047 -53
rect 1129 53 1175 100
rect 1129 19 1135 53
rect 1169 19 1175 53
rect 1129 -19 1175 19
rect 1129 -53 1135 -19
rect 1169 -53 1175 -19
rect 1129 -100 1175 -53
rect 1257 53 1303 100
rect 1257 19 1263 53
rect 1297 19 1303 53
rect 1257 -19 1303 19
rect 1257 -53 1263 -19
rect 1297 -53 1303 -19
rect 1257 -100 1303 -53
rect 1385 53 1431 100
rect 1385 19 1391 53
rect 1425 19 1431 53
rect 1385 -19 1431 19
rect 1385 -53 1391 -19
rect 1425 -53 1431 -19
rect 1385 -100 1431 -53
rect 1513 53 1559 100
rect 1513 19 1519 53
rect 1553 19 1559 53
rect 1513 -19 1559 19
rect 1513 -53 1519 -19
rect 1553 -53 1559 -19
rect 1513 -100 1559 -53
rect 1641 53 1687 100
rect 1641 19 1647 53
rect 1681 19 1687 53
rect 1641 -19 1687 19
rect 1641 -53 1647 -19
rect 1681 -53 1687 -19
rect 1641 -100 1687 -53
rect 1769 53 1815 100
rect 1769 19 1775 53
rect 1809 19 1815 53
rect 1769 -19 1815 19
rect 1769 -53 1775 -19
rect 1809 -53 1815 -19
rect 1769 -100 1815 -53
rect 1897 53 1943 100
rect 1897 19 1903 53
rect 1937 19 1943 53
rect 1897 -19 1943 19
rect 1897 -53 1903 -19
rect 1937 -53 1943 -19
rect 1897 -100 1943 -53
rect -1887 -147 -1825 -141
rect -1887 -181 -1873 -147
rect -1839 -181 -1825 -147
rect -1887 -187 -1825 -181
rect -1759 -147 -1697 -141
rect -1759 -181 -1745 -147
rect -1711 -181 -1697 -147
rect -1759 -187 -1697 -181
rect -1631 -147 -1569 -141
rect -1631 -181 -1617 -147
rect -1583 -181 -1569 -147
rect -1631 -187 -1569 -181
rect -1503 -147 -1441 -141
rect -1503 -181 -1489 -147
rect -1455 -181 -1441 -147
rect -1503 -187 -1441 -181
rect -1375 -147 -1313 -141
rect -1375 -181 -1361 -147
rect -1327 -181 -1313 -147
rect -1375 -187 -1313 -181
rect -1247 -147 -1185 -141
rect -1247 -181 -1233 -147
rect -1199 -181 -1185 -147
rect -1247 -187 -1185 -181
rect -1119 -147 -1057 -141
rect -1119 -181 -1105 -147
rect -1071 -181 -1057 -147
rect -1119 -187 -1057 -181
rect -991 -147 -929 -141
rect -991 -181 -977 -147
rect -943 -181 -929 -147
rect -991 -187 -929 -181
rect -863 -147 -801 -141
rect -863 -181 -849 -147
rect -815 -181 -801 -147
rect -863 -187 -801 -181
rect -735 -147 -673 -141
rect -735 -181 -721 -147
rect -687 -181 -673 -147
rect -735 -187 -673 -181
rect -607 -147 -545 -141
rect -607 -181 -593 -147
rect -559 -181 -545 -147
rect -607 -187 -545 -181
rect -479 -147 -417 -141
rect -479 -181 -465 -147
rect -431 -181 -417 -147
rect -479 -187 -417 -181
rect -351 -147 -289 -141
rect -351 -181 -337 -147
rect -303 -181 -289 -147
rect -351 -187 -289 -181
rect -223 -147 -161 -141
rect -223 -181 -209 -147
rect -175 -181 -161 -147
rect -223 -187 -161 -181
rect -95 -147 -33 -141
rect -95 -181 -81 -147
rect -47 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 47 -147
rect 81 -181 95 -147
rect 33 -187 95 -181
rect 161 -147 223 -141
rect 161 -181 175 -147
rect 209 -181 223 -147
rect 161 -187 223 -181
rect 289 -147 351 -141
rect 289 -181 303 -147
rect 337 -181 351 -147
rect 289 -187 351 -181
rect 417 -147 479 -141
rect 417 -181 431 -147
rect 465 -181 479 -147
rect 417 -187 479 -181
rect 545 -147 607 -141
rect 545 -181 559 -147
rect 593 -181 607 -147
rect 545 -187 607 -181
rect 673 -147 735 -141
rect 673 -181 687 -147
rect 721 -181 735 -147
rect 673 -187 735 -181
rect 801 -147 863 -141
rect 801 -181 815 -147
rect 849 -181 863 -147
rect 801 -187 863 -181
rect 929 -147 991 -141
rect 929 -181 943 -147
rect 977 -181 991 -147
rect 929 -187 991 -181
rect 1057 -147 1119 -141
rect 1057 -181 1071 -147
rect 1105 -181 1119 -147
rect 1057 -187 1119 -181
rect 1185 -147 1247 -141
rect 1185 -181 1199 -147
rect 1233 -181 1247 -147
rect 1185 -187 1247 -181
rect 1313 -147 1375 -141
rect 1313 -181 1327 -147
rect 1361 -181 1375 -147
rect 1313 -187 1375 -181
rect 1441 -147 1503 -141
rect 1441 -181 1455 -147
rect 1489 -181 1503 -147
rect 1441 -187 1503 -181
rect 1569 -147 1631 -141
rect 1569 -181 1583 -147
rect 1617 -181 1631 -147
rect 1569 -187 1631 -181
rect 1697 -147 1759 -141
rect 1697 -181 1711 -147
rect 1745 -181 1759 -147
rect 1697 -187 1759 -181
rect 1825 -147 1887 -141
rect 1825 -181 1839 -147
rect 1873 -181 1887 -147
rect 1825 -187 1887 -181
<< properties >>
string FIXED_BBOX -2034 -266 2034 266
<< end >>
