magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -3213 11102 3213 11188
rect -3213 -11102 -3127 11102
rect 3127 -11102 3213 11102
rect -3213 -11188 3213 -11102
<< psubdiff >>
rect -3187 11128 -3077 11162
rect -3043 11128 -3009 11162
rect -2975 11128 -2941 11162
rect -2907 11128 -2873 11162
rect -2839 11128 -2805 11162
rect -2771 11128 -2737 11162
rect -2703 11128 -2669 11162
rect -2635 11128 -2601 11162
rect -2567 11128 -2533 11162
rect -2499 11128 -2465 11162
rect -2431 11128 -2397 11162
rect -2363 11128 -2329 11162
rect -2295 11128 -2261 11162
rect -2227 11128 -2193 11162
rect -2159 11128 -2125 11162
rect -2091 11128 -2057 11162
rect -2023 11128 -1989 11162
rect -1955 11128 -1921 11162
rect -1887 11128 -1853 11162
rect -1819 11128 -1785 11162
rect -1751 11128 -1717 11162
rect -1683 11128 -1649 11162
rect -1615 11128 -1581 11162
rect -1547 11128 -1513 11162
rect -1479 11128 -1445 11162
rect -1411 11128 -1377 11162
rect -1343 11128 -1309 11162
rect -1275 11128 -1241 11162
rect -1207 11128 -1173 11162
rect -1139 11128 -1105 11162
rect -1071 11128 -1037 11162
rect -1003 11128 -969 11162
rect -935 11128 -901 11162
rect -867 11128 -833 11162
rect -799 11128 -765 11162
rect -731 11128 -697 11162
rect -663 11128 -629 11162
rect -595 11128 -561 11162
rect -527 11128 -493 11162
rect -459 11128 -425 11162
rect -391 11128 -357 11162
rect -323 11128 -289 11162
rect -255 11128 -221 11162
rect -187 11128 -153 11162
rect -119 11128 -85 11162
rect -51 11128 -17 11162
rect 17 11128 51 11162
rect 85 11128 119 11162
rect 153 11128 187 11162
rect 221 11128 255 11162
rect 289 11128 323 11162
rect 357 11128 391 11162
rect 425 11128 459 11162
rect 493 11128 527 11162
rect 561 11128 595 11162
rect 629 11128 663 11162
rect 697 11128 731 11162
rect 765 11128 799 11162
rect 833 11128 867 11162
rect 901 11128 935 11162
rect 969 11128 1003 11162
rect 1037 11128 1071 11162
rect 1105 11128 1139 11162
rect 1173 11128 1207 11162
rect 1241 11128 1275 11162
rect 1309 11128 1343 11162
rect 1377 11128 1411 11162
rect 1445 11128 1479 11162
rect 1513 11128 1547 11162
rect 1581 11128 1615 11162
rect 1649 11128 1683 11162
rect 1717 11128 1751 11162
rect 1785 11128 1819 11162
rect 1853 11128 1887 11162
rect 1921 11128 1955 11162
rect 1989 11128 2023 11162
rect 2057 11128 2091 11162
rect 2125 11128 2159 11162
rect 2193 11128 2227 11162
rect 2261 11128 2295 11162
rect 2329 11128 2363 11162
rect 2397 11128 2431 11162
rect 2465 11128 2499 11162
rect 2533 11128 2567 11162
rect 2601 11128 2635 11162
rect 2669 11128 2703 11162
rect 2737 11128 2771 11162
rect 2805 11128 2839 11162
rect 2873 11128 2907 11162
rect 2941 11128 2975 11162
rect 3009 11128 3043 11162
rect 3077 11128 3187 11162
rect -3187 11033 -3153 11128
rect 3153 11033 3187 11128
rect -3187 10965 -3153 10999
rect -3187 10897 -3153 10931
rect -3187 10829 -3153 10863
rect -3187 10761 -3153 10795
rect -3187 10693 -3153 10727
rect -3187 10625 -3153 10659
rect -3187 10557 -3153 10591
rect -3187 10489 -3153 10523
rect -3187 10421 -3153 10455
rect -3187 10353 -3153 10387
rect -3187 10285 -3153 10319
rect -3187 10217 -3153 10251
rect -3187 10149 -3153 10183
rect -3187 10081 -3153 10115
rect -3187 10013 -3153 10047
rect -3187 9945 -3153 9979
rect -3187 9877 -3153 9911
rect -3187 9809 -3153 9843
rect -3187 9741 -3153 9775
rect -3187 9673 -3153 9707
rect -3187 9605 -3153 9639
rect -3187 9537 -3153 9571
rect -3187 9469 -3153 9503
rect -3187 9401 -3153 9435
rect -3187 9333 -3153 9367
rect -3187 9265 -3153 9299
rect -3187 9197 -3153 9231
rect -3187 9129 -3153 9163
rect -3187 9061 -3153 9095
rect -3187 8993 -3153 9027
rect -3187 8925 -3153 8959
rect -3187 8857 -3153 8891
rect -3187 8789 -3153 8823
rect -3187 8721 -3153 8755
rect -3187 8653 -3153 8687
rect -3187 8585 -3153 8619
rect -3187 8517 -3153 8551
rect -3187 8449 -3153 8483
rect -3187 8381 -3153 8415
rect -3187 8313 -3153 8347
rect -3187 8245 -3153 8279
rect -3187 8177 -3153 8211
rect -3187 8109 -3153 8143
rect -3187 8041 -3153 8075
rect -3187 7973 -3153 8007
rect -3187 7905 -3153 7939
rect -3187 7837 -3153 7871
rect -3187 7769 -3153 7803
rect -3187 7701 -3153 7735
rect -3187 7633 -3153 7667
rect -3187 7565 -3153 7599
rect -3187 7497 -3153 7531
rect -3187 7429 -3153 7463
rect -3187 7361 -3153 7395
rect -3187 7293 -3153 7327
rect -3187 7225 -3153 7259
rect -3187 7157 -3153 7191
rect -3187 7089 -3153 7123
rect -3187 7021 -3153 7055
rect -3187 6953 -3153 6987
rect -3187 6885 -3153 6919
rect -3187 6817 -3153 6851
rect -3187 6749 -3153 6783
rect -3187 6681 -3153 6715
rect -3187 6613 -3153 6647
rect -3187 6545 -3153 6579
rect -3187 6477 -3153 6511
rect -3187 6409 -3153 6443
rect -3187 6341 -3153 6375
rect -3187 6273 -3153 6307
rect -3187 6205 -3153 6239
rect -3187 6137 -3153 6171
rect -3187 6069 -3153 6103
rect -3187 6001 -3153 6035
rect -3187 5933 -3153 5967
rect -3187 5865 -3153 5899
rect -3187 5797 -3153 5831
rect -3187 5729 -3153 5763
rect -3187 5661 -3153 5695
rect -3187 5593 -3153 5627
rect -3187 5525 -3153 5559
rect -3187 5457 -3153 5491
rect -3187 5389 -3153 5423
rect -3187 5321 -3153 5355
rect -3187 5253 -3153 5287
rect -3187 5185 -3153 5219
rect -3187 5117 -3153 5151
rect -3187 5049 -3153 5083
rect -3187 4981 -3153 5015
rect -3187 4913 -3153 4947
rect -3187 4845 -3153 4879
rect -3187 4777 -3153 4811
rect -3187 4709 -3153 4743
rect -3187 4641 -3153 4675
rect -3187 4573 -3153 4607
rect -3187 4505 -3153 4539
rect -3187 4437 -3153 4471
rect -3187 4369 -3153 4403
rect -3187 4301 -3153 4335
rect -3187 4233 -3153 4267
rect -3187 4165 -3153 4199
rect -3187 4097 -3153 4131
rect -3187 4029 -3153 4063
rect -3187 3961 -3153 3995
rect -3187 3893 -3153 3927
rect -3187 3825 -3153 3859
rect -3187 3757 -3153 3791
rect -3187 3689 -3153 3723
rect -3187 3621 -3153 3655
rect -3187 3553 -3153 3587
rect -3187 3485 -3153 3519
rect -3187 3417 -3153 3451
rect -3187 3349 -3153 3383
rect -3187 3281 -3153 3315
rect -3187 3213 -3153 3247
rect -3187 3145 -3153 3179
rect -3187 3077 -3153 3111
rect -3187 3009 -3153 3043
rect -3187 2941 -3153 2975
rect -3187 2873 -3153 2907
rect -3187 2805 -3153 2839
rect -3187 2737 -3153 2771
rect -3187 2669 -3153 2703
rect -3187 2601 -3153 2635
rect -3187 2533 -3153 2567
rect -3187 2465 -3153 2499
rect -3187 2397 -3153 2431
rect -3187 2329 -3153 2363
rect -3187 2261 -3153 2295
rect -3187 2193 -3153 2227
rect -3187 2125 -3153 2159
rect -3187 2057 -3153 2091
rect -3187 1989 -3153 2023
rect -3187 1921 -3153 1955
rect -3187 1853 -3153 1887
rect -3187 1785 -3153 1819
rect -3187 1717 -3153 1751
rect -3187 1649 -3153 1683
rect -3187 1581 -3153 1615
rect -3187 1513 -3153 1547
rect -3187 1445 -3153 1479
rect -3187 1377 -3153 1411
rect -3187 1309 -3153 1343
rect -3187 1241 -3153 1275
rect -3187 1173 -3153 1207
rect -3187 1105 -3153 1139
rect -3187 1037 -3153 1071
rect -3187 969 -3153 1003
rect -3187 901 -3153 935
rect -3187 833 -3153 867
rect -3187 765 -3153 799
rect -3187 697 -3153 731
rect -3187 629 -3153 663
rect -3187 561 -3153 595
rect -3187 493 -3153 527
rect -3187 425 -3153 459
rect -3187 357 -3153 391
rect -3187 289 -3153 323
rect -3187 221 -3153 255
rect -3187 153 -3153 187
rect -3187 85 -3153 119
rect -3187 17 -3153 51
rect -3187 -51 -3153 -17
rect -3187 -119 -3153 -85
rect -3187 -187 -3153 -153
rect -3187 -255 -3153 -221
rect -3187 -323 -3153 -289
rect -3187 -391 -3153 -357
rect -3187 -459 -3153 -425
rect -3187 -527 -3153 -493
rect -3187 -595 -3153 -561
rect -3187 -663 -3153 -629
rect -3187 -731 -3153 -697
rect -3187 -799 -3153 -765
rect -3187 -867 -3153 -833
rect -3187 -935 -3153 -901
rect -3187 -1003 -3153 -969
rect -3187 -1071 -3153 -1037
rect -3187 -1139 -3153 -1105
rect -3187 -1207 -3153 -1173
rect -3187 -1275 -3153 -1241
rect -3187 -1343 -3153 -1309
rect -3187 -1411 -3153 -1377
rect -3187 -1479 -3153 -1445
rect -3187 -1547 -3153 -1513
rect -3187 -1615 -3153 -1581
rect -3187 -1683 -3153 -1649
rect -3187 -1751 -3153 -1717
rect -3187 -1819 -3153 -1785
rect -3187 -1887 -3153 -1853
rect -3187 -1955 -3153 -1921
rect -3187 -2023 -3153 -1989
rect -3187 -2091 -3153 -2057
rect -3187 -2159 -3153 -2125
rect -3187 -2227 -3153 -2193
rect -3187 -2295 -3153 -2261
rect -3187 -2363 -3153 -2329
rect -3187 -2431 -3153 -2397
rect -3187 -2499 -3153 -2465
rect -3187 -2567 -3153 -2533
rect -3187 -2635 -3153 -2601
rect -3187 -2703 -3153 -2669
rect -3187 -2771 -3153 -2737
rect -3187 -2839 -3153 -2805
rect -3187 -2907 -3153 -2873
rect -3187 -2975 -3153 -2941
rect -3187 -3043 -3153 -3009
rect -3187 -3111 -3153 -3077
rect -3187 -3179 -3153 -3145
rect -3187 -3247 -3153 -3213
rect -3187 -3315 -3153 -3281
rect -3187 -3383 -3153 -3349
rect -3187 -3451 -3153 -3417
rect -3187 -3519 -3153 -3485
rect -3187 -3587 -3153 -3553
rect -3187 -3655 -3153 -3621
rect -3187 -3723 -3153 -3689
rect -3187 -3791 -3153 -3757
rect -3187 -3859 -3153 -3825
rect -3187 -3927 -3153 -3893
rect -3187 -3995 -3153 -3961
rect -3187 -4063 -3153 -4029
rect -3187 -4131 -3153 -4097
rect -3187 -4199 -3153 -4165
rect -3187 -4267 -3153 -4233
rect -3187 -4335 -3153 -4301
rect -3187 -4403 -3153 -4369
rect -3187 -4471 -3153 -4437
rect -3187 -4539 -3153 -4505
rect -3187 -4607 -3153 -4573
rect -3187 -4675 -3153 -4641
rect -3187 -4743 -3153 -4709
rect -3187 -4811 -3153 -4777
rect -3187 -4879 -3153 -4845
rect -3187 -4947 -3153 -4913
rect -3187 -5015 -3153 -4981
rect -3187 -5083 -3153 -5049
rect -3187 -5151 -3153 -5117
rect -3187 -5219 -3153 -5185
rect -3187 -5287 -3153 -5253
rect -3187 -5355 -3153 -5321
rect -3187 -5423 -3153 -5389
rect -3187 -5491 -3153 -5457
rect -3187 -5559 -3153 -5525
rect -3187 -5627 -3153 -5593
rect -3187 -5695 -3153 -5661
rect -3187 -5763 -3153 -5729
rect -3187 -5831 -3153 -5797
rect -3187 -5899 -3153 -5865
rect -3187 -5967 -3153 -5933
rect -3187 -6035 -3153 -6001
rect -3187 -6103 -3153 -6069
rect -3187 -6171 -3153 -6137
rect -3187 -6239 -3153 -6205
rect -3187 -6307 -3153 -6273
rect -3187 -6375 -3153 -6341
rect -3187 -6443 -3153 -6409
rect -3187 -6511 -3153 -6477
rect -3187 -6579 -3153 -6545
rect -3187 -6647 -3153 -6613
rect -3187 -6715 -3153 -6681
rect -3187 -6783 -3153 -6749
rect -3187 -6851 -3153 -6817
rect -3187 -6919 -3153 -6885
rect -3187 -6987 -3153 -6953
rect -3187 -7055 -3153 -7021
rect -3187 -7123 -3153 -7089
rect -3187 -7191 -3153 -7157
rect -3187 -7259 -3153 -7225
rect -3187 -7327 -3153 -7293
rect -3187 -7395 -3153 -7361
rect -3187 -7463 -3153 -7429
rect -3187 -7531 -3153 -7497
rect -3187 -7599 -3153 -7565
rect -3187 -7667 -3153 -7633
rect -3187 -7735 -3153 -7701
rect -3187 -7803 -3153 -7769
rect -3187 -7871 -3153 -7837
rect -3187 -7939 -3153 -7905
rect -3187 -8007 -3153 -7973
rect -3187 -8075 -3153 -8041
rect -3187 -8143 -3153 -8109
rect -3187 -8211 -3153 -8177
rect -3187 -8279 -3153 -8245
rect -3187 -8347 -3153 -8313
rect -3187 -8415 -3153 -8381
rect -3187 -8483 -3153 -8449
rect -3187 -8551 -3153 -8517
rect -3187 -8619 -3153 -8585
rect -3187 -8687 -3153 -8653
rect -3187 -8755 -3153 -8721
rect -3187 -8823 -3153 -8789
rect -3187 -8891 -3153 -8857
rect -3187 -8959 -3153 -8925
rect -3187 -9027 -3153 -8993
rect -3187 -9095 -3153 -9061
rect -3187 -9163 -3153 -9129
rect -3187 -9231 -3153 -9197
rect -3187 -9299 -3153 -9265
rect -3187 -9367 -3153 -9333
rect -3187 -9435 -3153 -9401
rect -3187 -9503 -3153 -9469
rect -3187 -9571 -3153 -9537
rect -3187 -9639 -3153 -9605
rect -3187 -9707 -3153 -9673
rect -3187 -9775 -3153 -9741
rect -3187 -9843 -3153 -9809
rect -3187 -9911 -3153 -9877
rect -3187 -9979 -3153 -9945
rect -3187 -10047 -3153 -10013
rect -3187 -10115 -3153 -10081
rect -3187 -10183 -3153 -10149
rect -3187 -10251 -3153 -10217
rect -3187 -10319 -3153 -10285
rect -3187 -10387 -3153 -10353
rect -3187 -10455 -3153 -10421
rect -3187 -10523 -3153 -10489
rect -3187 -10591 -3153 -10557
rect -3187 -10659 -3153 -10625
rect -3187 -10727 -3153 -10693
rect -3187 -10795 -3153 -10761
rect -3187 -10863 -3153 -10829
rect -3187 -10931 -3153 -10897
rect -3187 -10999 -3153 -10965
rect 3153 10965 3187 10999
rect 3153 10897 3187 10931
rect 3153 10829 3187 10863
rect 3153 10761 3187 10795
rect 3153 10693 3187 10727
rect 3153 10625 3187 10659
rect 3153 10557 3187 10591
rect 3153 10489 3187 10523
rect 3153 10421 3187 10455
rect 3153 10353 3187 10387
rect 3153 10285 3187 10319
rect 3153 10217 3187 10251
rect 3153 10149 3187 10183
rect 3153 10081 3187 10115
rect 3153 10013 3187 10047
rect 3153 9945 3187 9979
rect 3153 9877 3187 9911
rect 3153 9809 3187 9843
rect 3153 9741 3187 9775
rect 3153 9673 3187 9707
rect 3153 9605 3187 9639
rect 3153 9537 3187 9571
rect 3153 9469 3187 9503
rect 3153 9401 3187 9435
rect 3153 9333 3187 9367
rect 3153 9265 3187 9299
rect 3153 9197 3187 9231
rect 3153 9129 3187 9163
rect 3153 9061 3187 9095
rect 3153 8993 3187 9027
rect 3153 8925 3187 8959
rect 3153 8857 3187 8891
rect 3153 8789 3187 8823
rect 3153 8721 3187 8755
rect 3153 8653 3187 8687
rect 3153 8585 3187 8619
rect 3153 8517 3187 8551
rect 3153 8449 3187 8483
rect 3153 8381 3187 8415
rect 3153 8313 3187 8347
rect 3153 8245 3187 8279
rect 3153 8177 3187 8211
rect 3153 8109 3187 8143
rect 3153 8041 3187 8075
rect 3153 7973 3187 8007
rect 3153 7905 3187 7939
rect 3153 7837 3187 7871
rect 3153 7769 3187 7803
rect 3153 7701 3187 7735
rect 3153 7633 3187 7667
rect 3153 7565 3187 7599
rect 3153 7497 3187 7531
rect 3153 7429 3187 7463
rect 3153 7361 3187 7395
rect 3153 7293 3187 7327
rect 3153 7225 3187 7259
rect 3153 7157 3187 7191
rect 3153 7089 3187 7123
rect 3153 7021 3187 7055
rect 3153 6953 3187 6987
rect 3153 6885 3187 6919
rect 3153 6817 3187 6851
rect 3153 6749 3187 6783
rect 3153 6681 3187 6715
rect 3153 6613 3187 6647
rect 3153 6545 3187 6579
rect 3153 6477 3187 6511
rect 3153 6409 3187 6443
rect 3153 6341 3187 6375
rect 3153 6273 3187 6307
rect 3153 6205 3187 6239
rect 3153 6137 3187 6171
rect 3153 6069 3187 6103
rect 3153 6001 3187 6035
rect 3153 5933 3187 5967
rect 3153 5865 3187 5899
rect 3153 5797 3187 5831
rect 3153 5729 3187 5763
rect 3153 5661 3187 5695
rect 3153 5593 3187 5627
rect 3153 5525 3187 5559
rect 3153 5457 3187 5491
rect 3153 5389 3187 5423
rect 3153 5321 3187 5355
rect 3153 5253 3187 5287
rect 3153 5185 3187 5219
rect 3153 5117 3187 5151
rect 3153 5049 3187 5083
rect 3153 4981 3187 5015
rect 3153 4913 3187 4947
rect 3153 4845 3187 4879
rect 3153 4777 3187 4811
rect 3153 4709 3187 4743
rect 3153 4641 3187 4675
rect 3153 4573 3187 4607
rect 3153 4505 3187 4539
rect 3153 4437 3187 4471
rect 3153 4369 3187 4403
rect 3153 4301 3187 4335
rect 3153 4233 3187 4267
rect 3153 4165 3187 4199
rect 3153 4097 3187 4131
rect 3153 4029 3187 4063
rect 3153 3961 3187 3995
rect 3153 3893 3187 3927
rect 3153 3825 3187 3859
rect 3153 3757 3187 3791
rect 3153 3689 3187 3723
rect 3153 3621 3187 3655
rect 3153 3553 3187 3587
rect 3153 3485 3187 3519
rect 3153 3417 3187 3451
rect 3153 3349 3187 3383
rect 3153 3281 3187 3315
rect 3153 3213 3187 3247
rect 3153 3145 3187 3179
rect 3153 3077 3187 3111
rect 3153 3009 3187 3043
rect 3153 2941 3187 2975
rect 3153 2873 3187 2907
rect 3153 2805 3187 2839
rect 3153 2737 3187 2771
rect 3153 2669 3187 2703
rect 3153 2601 3187 2635
rect 3153 2533 3187 2567
rect 3153 2465 3187 2499
rect 3153 2397 3187 2431
rect 3153 2329 3187 2363
rect 3153 2261 3187 2295
rect 3153 2193 3187 2227
rect 3153 2125 3187 2159
rect 3153 2057 3187 2091
rect 3153 1989 3187 2023
rect 3153 1921 3187 1955
rect 3153 1853 3187 1887
rect 3153 1785 3187 1819
rect 3153 1717 3187 1751
rect 3153 1649 3187 1683
rect 3153 1581 3187 1615
rect 3153 1513 3187 1547
rect 3153 1445 3187 1479
rect 3153 1377 3187 1411
rect 3153 1309 3187 1343
rect 3153 1241 3187 1275
rect 3153 1173 3187 1207
rect 3153 1105 3187 1139
rect 3153 1037 3187 1071
rect 3153 969 3187 1003
rect 3153 901 3187 935
rect 3153 833 3187 867
rect 3153 765 3187 799
rect 3153 697 3187 731
rect 3153 629 3187 663
rect 3153 561 3187 595
rect 3153 493 3187 527
rect 3153 425 3187 459
rect 3153 357 3187 391
rect 3153 289 3187 323
rect 3153 221 3187 255
rect 3153 153 3187 187
rect 3153 85 3187 119
rect 3153 17 3187 51
rect 3153 -51 3187 -17
rect 3153 -119 3187 -85
rect 3153 -187 3187 -153
rect 3153 -255 3187 -221
rect 3153 -323 3187 -289
rect 3153 -391 3187 -357
rect 3153 -459 3187 -425
rect 3153 -527 3187 -493
rect 3153 -595 3187 -561
rect 3153 -663 3187 -629
rect 3153 -731 3187 -697
rect 3153 -799 3187 -765
rect 3153 -867 3187 -833
rect 3153 -935 3187 -901
rect 3153 -1003 3187 -969
rect 3153 -1071 3187 -1037
rect 3153 -1139 3187 -1105
rect 3153 -1207 3187 -1173
rect 3153 -1275 3187 -1241
rect 3153 -1343 3187 -1309
rect 3153 -1411 3187 -1377
rect 3153 -1479 3187 -1445
rect 3153 -1547 3187 -1513
rect 3153 -1615 3187 -1581
rect 3153 -1683 3187 -1649
rect 3153 -1751 3187 -1717
rect 3153 -1819 3187 -1785
rect 3153 -1887 3187 -1853
rect 3153 -1955 3187 -1921
rect 3153 -2023 3187 -1989
rect 3153 -2091 3187 -2057
rect 3153 -2159 3187 -2125
rect 3153 -2227 3187 -2193
rect 3153 -2295 3187 -2261
rect 3153 -2363 3187 -2329
rect 3153 -2431 3187 -2397
rect 3153 -2499 3187 -2465
rect 3153 -2567 3187 -2533
rect 3153 -2635 3187 -2601
rect 3153 -2703 3187 -2669
rect 3153 -2771 3187 -2737
rect 3153 -2839 3187 -2805
rect 3153 -2907 3187 -2873
rect 3153 -2975 3187 -2941
rect 3153 -3043 3187 -3009
rect 3153 -3111 3187 -3077
rect 3153 -3179 3187 -3145
rect 3153 -3247 3187 -3213
rect 3153 -3315 3187 -3281
rect 3153 -3383 3187 -3349
rect 3153 -3451 3187 -3417
rect 3153 -3519 3187 -3485
rect 3153 -3587 3187 -3553
rect 3153 -3655 3187 -3621
rect 3153 -3723 3187 -3689
rect 3153 -3791 3187 -3757
rect 3153 -3859 3187 -3825
rect 3153 -3927 3187 -3893
rect 3153 -3995 3187 -3961
rect 3153 -4063 3187 -4029
rect 3153 -4131 3187 -4097
rect 3153 -4199 3187 -4165
rect 3153 -4267 3187 -4233
rect 3153 -4335 3187 -4301
rect 3153 -4403 3187 -4369
rect 3153 -4471 3187 -4437
rect 3153 -4539 3187 -4505
rect 3153 -4607 3187 -4573
rect 3153 -4675 3187 -4641
rect 3153 -4743 3187 -4709
rect 3153 -4811 3187 -4777
rect 3153 -4879 3187 -4845
rect 3153 -4947 3187 -4913
rect 3153 -5015 3187 -4981
rect 3153 -5083 3187 -5049
rect 3153 -5151 3187 -5117
rect 3153 -5219 3187 -5185
rect 3153 -5287 3187 -5253
rect 3153 -5355 3187 -5321
rect 3153 -5423 3187 -5389
rect 3153 -5491 3187 -5457
rect 3153 -5559 3187 -5525
rect 3153 -5627 3187 -5593
rect 3153 -5695 3187 -5661
rect 3153 -5763 3187 -5729
rect 3153 -5831 3187 -5797
rect 3153 -5899 3187 -5865
rect 3153 -5967 3187 -5933
rect 3153 -6035 3187 -6001
rect 3153 -6103 3187 -6069
rect 3153 -6171 3187 -6137
rect 3153 -6239 3187 -6205
rect 3153 -6307 3187 -6273
rect 3153 -6375 3187 -6341
rect 3153 -6443 3187 -6409
rect 3153 -6511 3187 -6477
rect 3153 -6579 3187 -6545
rect 3153 -6647 3187 -6613
rect 3153 -6715 3187 -6681
rect 3153 -6783 3187 -6749
rect 3153 -6851 3187 -6817
rect 3153 -6919 3187 -6885
rect 3153 -6987 3187 -6953
rect 3153 -7055 3187 -7021
rect 3153 -7123 3187 -7089
rect 3153 -7191 3187 -7157
rect 3153 -7259 3187 -7225
rect 3153 -7327 3187 -7293
rect 3153 -7395 3187 -7361
rect 3153 -7463 3187 -7429
rect 3153 -7531 3187 -7497
rect 3153 -7599 3187 -7565
rect 3153 -7667 3187 -7633
rect 3153 -7735 3187 -7701
rect 3153 -7803 3187 -7769
rect 3153 -7871 3187 -7837
rect 3153 -7939 3187 -7905
rect 3153 -8007 3187 -7973
rect 3153 -8075 3187 -8041
rect 3153 -8143 3187 -8109
rect 3153 -8211 3187 -8177
rect 3153 -8279 3187 -8245
rect 3153 -8347 3187 -8313
rect 3153 -8415 3187 -8381
rect 3153 -8483 3187 -8449
rect 3153 -8551 3187 -8517
rect 3153 -8619 3187 -8585
rect 3153 -8687 3187 -8653
rect 3153 -8755 3187 -8721
rect 3153 -8823 3187 -8789
rect 3153 -8891 3187 -8857
rect 3153 -8959 3187 -8925
rect 3153 -9027 3187 -8993
rect 3153 -9095 3187 -9061
rect 3153 -9163 3187 -9129
rect 3153 -9231 3187 -9197
rect 3153 -9299 3187 -9265
rect 3153 -9367 3187 -9333
rect 3153 -9435 3187 -9401
rect 3153 -9503 3187 -9469
rect 3153 -9571 3187 -9537
rect 3153 -9639 3187 -9605
rect 3153 -9707 3187 -9673
rect 3153 -9775 3187 -9741
rect 3153 -9843 3187 -9809
rect 3153 -9911 3187 -9877
rect 3153 -9979 3187 -9945
rect 3153 -10047 3187 -10013
rect 3153 -10115 3187 -10081
rect 3153 -10183 3187 -10149
rect 3153 -10251 3187 -10217
rect 3153 -10319 3187 -10285
rect 3153 -10387 3187 -10353
rect 3153 -10455 3187 -10421
rect 3153 -10523 3187 -10489
rect 3153 -10591 3187 -10557
rect 3153 -10659 3187 -10625
rect 3153 -10727 3187 -10693
rect 3153 -10795 3187 -10761
rect 3153 -10863 3187 -10829
rect 3153 -10931 3187 -10897
rect 3153 -10999 3187 -10965
rect -3187 -11128 -3153 -11033
rect 3153 -11128 3187 -11033
rect -3187 -11162 -3077 -11128
rect -3043 -11162 -3009 -11128
rect -2975 -11162 -2941 -11128
rect -2907 -11162 -2873 -11128
rect -2839 -11162 -2805 -11128
rect -2771 -11162 -2737 -11128
rect -2703 -11162 -2669 -11128
rect -2635 -11162 -2601 -11128
rect -2567 -11162 -2533 -11128
rect -2499 -11162 -2465 -11128
rect -2431 -11162 -2397 -11128
rect -2363 -11162 -2329 -11128
rect -2295 -11162 -2261 -11128
rect -2227 -11162 -2193 -11128
rect -2159 -11162 -2125 -11128
rect -2091 -11162 -2057 -11128
rect -2023 -11162 -1989 -11128
rect -1955 -11162 -1921 -11128
rect -1887 -11162 -1853 -11128
rect -1819 -11162 -1785 -11128
rect -1751 -11162 -1717 -11128
rect -1683 -11162 -1649 -11128
rect -1615 -11162 -1581 -11128
rect -1547 -11162 -1513 -11128
rect -1479 -11162 -1445 -11128
rect -1411 -11162 -1377 -11128
rect -1343 -11162 -1309 -11128
rect -1275 -11162 -1241 -11128
rect -1207 -11162 -1173 -11128
rect -1139 -11162 -1105 -11128
rect -1071 -11162 -1037 -11128
rect -1003 -11162 -969 -11128
rect -935 -11162 -901 -11128
rect -867 -11162 -833 -11128
rect -799 -11162 -765 -11128
rect -731 -11162 -697 -11128
rect -663 -11162 -629 -11128
rect -595 -11162 -561 -11128
rect -527 -11162 -493 -11128
rect -459 -11162 -425 -11128
rect -391 -11162 -357 -11128
rect -323 -11162 -289 -11128
rect -255 -11162 -221 -11128
rect -187 -11162 -153 -11128
rect -119 -11162 -85 -11128
rect -51 -11162 -17 -11128
rect 17 -11162 51 -11128
rect 85 -11162 119 -11128
rect 153 -11162 187 -11128
rect 221 -11162 255 -11128
rect 289 -11162 323 -11128
rect 357 -11162 391 -11128
rect 425 -11162 459 -11128
rect 493 -11162 527 -11128
rect 561 -11162 595 -11128
rect 629 -11162 663 -11128
rect 697 -11162 731 -11128
rect 765 -11162 799 -11128
rect 833 -11162 867 -11128
rect 901 -11162 935 -11128
rect 969 -11162 1003 -11128
rect 1037 -11162 1071 -11128
rect 1105 -11162 1139 -11128
rect 1173 -11162 1207 -11128
rect 1241 -11162 1275 -11128
rect 1309 -11162 1343 -11128
rect 1377 -11162 1411 -11128
rect 1445 -11162 1479 -11128
rect 1513 -11162 1547 -11128
rect 1581 -11162 1615 -11128
rect 1649 -11162 1683 -11128
rect 1717 -11162 1751 -11128
rect 1785 -11162 1819 -11128
rect 1853 -11162 1887 -11128
rect 1921 -11162 1955 -11128
rect 1989 -11162 2023 -11128
rect 2057 -11162 2091 -11128
rect 2125 -11162 2159 -11128
rect 2193 -11162 2227 -11128
rect 2261 -11162 2295 -11128
rect 2329 -11162 2363 -11128
rect 2397 -11162 2431 -11128
rect 2465 -11162 2499 -11128
rect 2533 -11162 2567 -11128
rect 2601 -11162 2635 -11128
rect 2669 -11162 2703 -11128
rect 2737 -11162 2771 -11128
rect 2805 -11162 2839 -11128
rect 2873 -11162 2907 -11128
rect 2941 -11162 2975 -11128
rect 3009 -11162 3043 -11128
rect 3077 -11162 3187 -11128
<< psubdiffcont >>
rect -3077 11128 -3043 11162
rect -3009 11128 -2975 11162
rect -2941 11128 -2907 11162
rect -2873 11128 -2839 11162
rect -2805 11128 -2771 11162
rect -2737 11128 -2703 11162
rect -2669 11128 -2635 11162
rect -2601 11128 -2567 11162
rect -2533 11128 -2499 11162
rect -2465 11128 -2431 11162
rect -2397 11128 -2363 11162
rect -2329 11128 -2295 11162
rect -2261 11128 -2227 11162
rect -2193 11128 -2159 11162
rect -2125 11128 -2091 11162
rect -2057 11128 -2023 11162
rect -1989 11128 -1955 11162
rect -1921 11128 -1887 11162
rect -1853 11128 -1819 11162
rect -1785 11128 -1751 11162
rect -1717 11128 -1683 11162
rect -1649 11128 -1615 11162
rect -1581 11128 -1547 11162
rect -1513 11128 -1479 11162
rect -1445 11128 -1411 11162
rect -1377 11128 -1343 11162
rect -1309 11128 -1275 11162
rect -1241 11128 -1207 11162
rect -1173 11128 -1139 11162
rect -1105 11128 -1071 11162
rect -1037 11128 -1003 11162
rect -969 11128 -935 11162
rect -901 11128 -867 11162
rect -833 11128 -799 11162
rect -765 11128 -731 11162
rect -697 11128 -663 11162
rect -629 11128 -595 11162
rect -561 11128 -527 11162
rect -493 11128 -459 11162
rect -425 11128 -391 11162
rect -357 11128 -323 11162
rect -289 11128 -255 11162
rect -221 11128 -187 11162
rect -153 11128 -119 11162
rect -85 11128 -51 11162
rect -17 11128 17 11162
rect 51 11128 85 11162
rect 119 11128 153 11162
rect 187 11128 221 11162
rect 255 11128 289 11162
rect 323 11128 357 11162
rect 391 11128 425 11162
rect 459 11128 493 11162
rect 527 11128 561 11162
rect 595 11128 629 11162
rect 663 11128 697 11162
rect 731 11128 765 11162
rect 799 11128 833 11162
rect 867 11128 901 11162
rect 935 11128 969 11162
rect 1003 11128 1037 11162
rect 1071 11128 1105 11162
rect 1139 11128 1173 11162
rect 1207 11128 1241 11162
rect 1275 11128 1309 11162
rect 1343 11128 1377 11162
rect 1411 11128 1445 11162
rect 1479 11128 1513 11162
rect 1547 11128 1581 11162
rect 1615 11128 1649 11162
rect 1683 11128 1717 11162
rect 1751 11128 1785 11162
rect 1819 11128 1853 11162
rect 1887 11128 1921 11162
rect 1955 11128 1989 11162
rect 2023 11128 2057 11162
rect 2091 11128 2125 11162
rect 2159 11128 2193 11162
rect 2227 11128 2261 11162
rect 2295 11128 2329 11162
rect 2363 11128 2397 11162
rect 2431 11128 2465 11162
rect 2499 11128 2533 11162
rect 2567 11128 2601 11162
rect 2635 11128 2669 11162
rect 2703 11128 2737 11162
rect 2771 11128 2805 11162
rect 2839 11128 2873 11162
rect 2907 11128 2941 11162
rect 2975 11128 3009 11162
rect 3043 11128 3077 11162
rect -3187 10999 -3153 11033
rect -3187 10931 -3153 10965
rect -3187 10863 -3153 10897
rect -3187 10795 -3153 10829
rect -3187 10727 -3153 10761
rect -3187 10659 -3153 10693
rect -3187 10591 -3153 10625
rect -3187 10523 -3153 10557
rect -3187 10455 -3153 10489
rect -3187 10387 -3153 10421
rect -3187 10319 -3153 10353
rect -3187 10251 -3153 10285
rect -3187 10183 -3153 10217
rect -3187 10115 -3153 10149
rect -3187 10047 -3153 10081
rect -3187 9979 -3153 10013
rect -3187 9911 -3153 9945
rect -3187 9843 -3153 9877
rect -3187 9775 -3153 9809
rect -3187 9707 -3153 9741
rect -3187 9639 -3153 9673
rect -3187 9571 -3153 9605
rect -3187 9503 -3153 9537
rect -3187 9435 -3153 9469
rect -3187 9367 -3153 9401
rect -3187 9299 -3153 9333
rect -3187 9231 -3153 9265
rect -3187 9163 -3153 9197
rect -3187 9095 -3153 9129
rect -3187 9027 -3153 9061
rect -3187 8959 -3153 8993
rect -3187 8891 -3153 8925
rect -3187 8823 -3153 8857
rect -3187 8755 -3153 8789
rect -3187 8687 -3153 8721
rect -3187 8619 -3153 8653
rect -3187 8551 -3153 8585
rect -3187 8483 -3153 8517
rect -3187 8415 -3153 8449
rect -3187 8347 -3153 8381
rect -3187 8279 -3153 8313
rect -3187 8211 -3153 8245
rect -3187 8143 -3153 8177
rect -3187 8075 -3153 8109
rect -3187 8007 -3153 8041
rect -3187 7939 -3153 7973
rect -3187 7871 -3153 7905
rect -3187 7803 -3153 7837
rect -3187 7735 -3153 7769
rect -3187 7667 -3153 7701
rect -3187 7599 -3153 7633
rect -3187 7531 -3153 7565
rect -3187 7463 -3153 7497
rect -3187 7395 -3153 7429
rect -3187 7327 -3153 7361
rect -3187 7259 -3153 7293
rect -3187 7191 -3153 7225
rect -3187 7123 -3153 7157
rect -3187 7055 -3153 7089
rect -3187 6987 -3153 7021
rect -3187 6919 -3153 6953
rect -3187 6851 -3153 6885
rect -3187 6783 -3153 6817
rect -3187 6715 -3153 6749
rect -3187 6647 -3153 6681
rect -3187 6579 -3153 6613
rect -3187 6511 -3153 6545
rect -3187 6443 -3153 6477
rect -3187 6375 -3153 6409
rect -3187 6307 -3153 6341
rect -3187 6239 -3153 6273
rect -3187 6171 -3153 6205
rect -3187 6103 -3153 6137
rect -3187 6035 -3153 6069
rect -3187 5967 -3153 6001
rect -3187 5899 -3153 5933
rect -3187 5831 -3153 5865
rect -3187 5763 -3153 5797
rect -3187 5695 -3153 5729
rect -3187 5627 -3153 5661
rect -3187 5559 -3153 5593
rect -3187 5491 -3153 5525
rect -3187 5423 -3153 5457
rect -3187 5355 -3153 5389
rect -3187 5287 -3153 5321
rect -3187 5219 -3153 5253
rect -3187 5151 -3153 5185
rect -3187 5083 -3153 5117
rect -3187 5015 -3153 5049
rect -3187 4947 -3153 4981
rect -3187 4879 -3153 4913
rect -3187 4811 -3153 4845
rect -3187 4743 -3153 4777
rect -3187 4675 -3153 4709
rect -3187 4607 -3153 4641
rect -3187 4539 -3153 4573
rect -3187 4471 -3153 4505
rect -3187 4403 -3153 4437
rect -3187 4335 -3153 4369
rect -3187 4267 -3153 4301
rect -3187 4199 -3153 4233
rect -3187 4131 -3153 4165
rect -3187 4063 -3153 4097
rect -3187 3995 -3153 4029
rect -3187 3927 -3153 3961
rect -3187 3859 -3153 3893
rect -3187 3791 -3153 3825
rect -3187 3723 -3153 3757
rect -3187 3655 -3153 3689
rect -3187 3587 -3153 3621
rect -3187 3519 -3153 3553
rect -3187 3451 -3153 3485
rect -3187 3383 -3153 3417
rect -3187 3315 -3153 3349
rect -3187 3247 -3153 3281
rect -3187 3179 -3153 3213
rect -3187 3111 -3153 3145
rect -3187 3043 -3153 3077
rect -3187 2975 -3153 3009
rect -3187 2907 -3153 2941
rect -3187 2839 -3153 2873
rect -3187 2771 -3153 2805
rect -3187 2703 -3153 2737
rect -3187 2635 -3153 2669
rect -3187 2567 -3153 2601
rect -3187 2499 -3153 2533
rect -3187 2431 -3153 2465
rect -3187 2363 -3153 2397
rect -3187 2295 -3153 2329
rect -3187 2227 -3153 2261
rect -3187 2159 -3153 2193
rect -3187 2091 -3153 2125
rect -3187 2023 -3153 2057
rect -3187 1955 -3153 1989
rect -3187 1887 -3153 1921
rect -3187 1819 -3153 1853
rect -3187 1751 -3153 1785
rect -3187 1683 -3153 1717
rect -3187 1615 -3153 1649
rect -3187 1547 -3153 1581
rect -3187 1479 -3153 1513
rect -3187 1411 -3153 1445
rect -3187 1343 -3153 1377
rect -3187 1275 -3153 1309
rect -3187 1207 -3153 1241
rect -3187 1139 -3153 1173
rect -3187 1071 -3153 1105
rect -3187 1003 -3153 1037
rect -3187 935 -3153 969
rect -3187 867 -3153 901
rect -3187 799 -3153 833
rect -3187 731 -3153 765
rect -3187 663 -3153 697
rect -3187 595 -3153 629
rect -3187 527 -3153 561
rect -3187 459 -3153 493
rect -3187 391 -3153 425
rect -3187 323 -3153 357
rect -3187 255 -3153 289
rect -3187 187 -3153 221
rect -3187 119 -3153 153
rect -3187 51 -3153 85
rect -3187 -17 -3153 17
rect -3187 -85 -3153 -51
rect -3187 -153 -3153 -119
rect -3187 -221 -3153 -187
rect -3187 -289 -3153 -255
rect -3187 -357 -3153 -323
rect -3187 -425 -3153 -391
rect -3187 -493 -3153 -459
rect -3187 -561 -3153 -527
rect -3187 -629 -3153 -595
rect -3187 -697 -3153 -663
rect -3187 -765 -3153 -731
rect -3187 -833 -3153 -799
rect -3187 -901 -3153 -867
rect -3187 -969 -3153 -935
rect -3187 -1037 -3153 -1003
rect -3187 -1105 -3153 -1071
rect -3187 -1173 -3153 -1139
rect -3187 -1241 -3153 -1207
rect -3187 -1309 -3153 -1275
rect -3187 -1377 -3153 -1343
rect -3187 -1445 -3153 -1411
rect -3187 -1513 -3153 -1479
rect -3187 -1581 -3153 -1547
rect -3187 -1649 -3153 -1615
rect -3187 -1717 -3153 -1683
rect -3187 -1785 -3153 -1751
rect -3187 -1853 -3153 -1819
rect -3187 -1921 -3153 -1887
rect -3187 -1989 -3153 -1955
rect -3187 -2057 -3153 -2023
rect -3187 -2125 -3153 -2091
rect -3187 -2193 -3153 -2159
rect -3187 -2261 -3153 -2227
rect -3187 -2329 -3153 -2295
rect -3187 -2397 -3153 -2363
rect -3187 -2465 -3153 -2431
rect -3187 -2533 -3153 -2499
rect -3187 -2601 -3153 -2567
rect -3187 -2669 -3153 -2635
rect -3187 -2737 -3153 -2703
rect -3187 -2805 -3153 -2771
rect -3187 -2873 -3153 -2839
rect -3187 -2941 -3153 -2907
rect -3187 -3009 -3153 -2975
rect -3187 -3077 -3153 -3043
rect -3187 -3145 -3153 -3111
rect -3187 -3213 -3153 -3179
rect -3187 -3281 -3153 -3247
rect -3187 -3349 -3153 -3315
rect -3187 -3417 -3153 -3383
rect -3187 -3485 -3153 -3451
rect -3187 -3553 -3153 -3519
rect -3187 -3621 -3153 -3587
rect -3187 -3689 -3153 -3655
rect -3187 -3757 -3153 -3723
rect -3187 -3825 -3153 -3791
rect -3187 -3893 -3153 -3859
rect -3187 -3961 -3153 -3927
rect -3187 -4029 -3153 -3995
rect -3187 -4097 -3153 -4063
rect -3187 -4165 -3153 -4131
rect -3187 -4233 -3153 -4199
rect -3187 -4301 -3153 -4267
rect -3187 -4369 -3153 -4335
rect -3187 -4437 -3153 -4403
rect -3187 -4505 -3153 -4471
rect -3187 -4573 -3153 -4539
rect -3187 -4641 -3153 -4607
rect -3187 -4709 -3153 -4675
rect -3187 -4777 -3153 -4743
rect -3187 -4845 -3153 -4811
rect -3187 -4913 -3153 -4879
rect -3187 -4981 -3153 -4947
rect -3187 -5049 -3153 -5015
rect -3187 -5117 -3153 -5083
rect -3187 -5185 -3153 -5151
rect -3187 -5253 -3153 -5219
rect -3187 -5321 -3153 -5287
rect -3187 -5389 -3153 -5355
rect -3187 -5457 -3153 -5423
rect -3187 -5525 -3153 -5491
rect -3187 -5593 -3153 -5559
rect -3187 -5661 -3153 -5627
rect -3187 -5729 -3153 -5695
rect -3187 -5797 -3153 -5763
rect -3187 -5865 -3153 -5831
rect -3187 -5933 -3153 -5899
rect -3187 -6001 -3153 -5967
rect -3187 -6069 -3153 -6035
rect -3187 -6137 -3153 -6103
rect -3187 -6205 -3153 -6171
rect -3187 -6273 -3153 -6239
rect -3187 -6341 -3153 -6307
rect -3187 -6409 -3153 -6375
rect -3187 -6477 -3153 -6443
rect -3187 -6545 -3153 -6511
rect -3187 -6613 -3153 -6579
rect -3187 -6681 -3153 -6647
rect -3187 -6749 -3153 -6715
rect -3187 -6817 -3153 -6783
rect -3187 -6885 -3153 -6851
rect -3187 -6953 -3153 -6919
rect -3187 -7021 -3153 -6987
rect -3187 -7089 -3153 -7055
rect -3187 -7157 -3153 -7123
rect -3187 -7225 -3153 -7191
rect -3187 -7293 -3153 -7259
rect -3187 -7361 -3153 -7327
rect -3187 -7429 -3153 -7395
rect -3187 -7497 -3153 -7463
rect -3187 -7565 -3153 -7531
rect -3187 -7633 -3153 -7599
rect -3187 -7701 -3153 -7667
rect -3187 -7769 -3153 -7735
rect -3187 -7837 -3153 -7803
rect -3187 -7905 -3153 -7871
rect -3187 -7973 -3153 -7939
rect -3187 -8041 -3153 -8007
rect -3187 -8109 -3153 -8075
rect -3187 -8177 -3153 -8143
rect -3187 -8245 -3153 -8211
rect -3187 -8313 -3153 -8279
rect -3187 -8381 -3153 -8347
rect -3187 -8449 -3153 -8415
rect -3187 -8517 -3153 -8483
rect -3187 -8585 -3153 -8551
rect -3187 -8653 -3153 -8619
rect -3187 -8721 -3153 -8687
rect -3187 -8789 -3153 -8755
rect -3187 -8857 -3153 -8823
rect -3187 -8925 -3153 -8891
rect -3187 -8993 -3153 -8959
rect -3187 -9061 -3153 -9027
rect -3187 -9129 -3153 -9095
rect -3187 -9197 -3153 -9163
rect -3187 -9265 -3153 -9231
rect -3187 -9333 -3153 -9299
rect -3187 -9401 -3153 -9367
rect -3187 -9469 -3153 -9435
rect -3187 -9537 -3153 -9503
rect -3187 -9605 -3153 -9571
rect -3187 -9673 -3153 -9639
rect -3187 -9741 -3153 -9707
rect -3187 -9809 -3153 -9775
rect -3187 -9877 -3153 -9843
rect -3187 -9945 -3153 -9911
rect -3187 -10013 -3153 -9979
rect -3187 -10081 -3153 -10047
rect -3187 -10149 -3153 -10115
rect -3187 -10217 -3153 -10183
rect -3187 -10285 -3153 -10251
rect -3187 -10353 -3153 -10319
rect -3187 -10421 -3153 -10387
rect -3187 -10489 -3153 -10455
rect -3187 -10557 -3153 -10523
rect -3187 -10625 -3153 -10591
rect -3187 -10693 -3153 -10659
rect -3187 -10761 -3153 -10727
rect -3187 -10829 -3153 -10795
rect -3187 -10897 -3153 -10863
rect -3187 -10965 -3153 -10931
rect -3187 -11033 -3153 -10999
rect 3153 10999 3187 11033
rect 3153 10931 3187 10965
rect 3153 10863 3187 10897
rect 3153 10795 3187 10829
rect 3153 10727 3187 10761
rect 3153 10659 3187 10693
rect 3153 10591 3187 10625
rect 3153 10523 3187 10557
rect 3153 10455 3187 10489
rect 3153 10387 3187 10421
rect 3153 10319 3187 10353
rect 3153 10251 3187 10285
rect 3153 10183 3187 10217
rect 3153 10115 3187 10149
rect 3153 10047 3187 10081
rect 3153 9979 3187 10013
rect 3153 9911 3187 9945
rect 3153 9843 3187 9877
rect 3153 9775 3187 9809
rect 3153 9707 3187 9741
rect 3153 9639 3187 9673
rect 3153 9571 3187 9605
rect 3153 9503 3187 9537
rect 3153 9435 3187 9469
rect 3153 9367 3187 9401
rect 3153 9299 3187 9333
rect 3153 9231 3187 9265
rect 3153 9163 3187 9197
rect 3153 9095 3187 9129
rect 3153 9027 3187 9061
rect 3153 8959 3187 8993
rect 3153 8891 3187 8925
rect 3153 8823 3187 8857
rect 3153 8755 3187 8789
rect 3153 8687 3187 8721
rect 3153 8619 3187 8653
rect 3153 8551 3187 8585
rect 3153 8483 3187 8517
rect 3153 8415 3187 8449
rect 3153 8347 3187 8381
rect 3153 8279 3187 8313
rect 3153 8211 3187 8245
rect 3153 8143 3187 8177
rect 3153 8075 3187 8109
rect 3153 8007 3187 8041
rect 3153 7939 3187 7973
rect 3153 7871 3187 7905
rect 3153 7803 3187 7837
rect 3153 7735 3187 7769
rect 3153 7667 3187 7701
rect 3153 7599 3187 7633
rect 3153 7531 3187 7565
rect 3153 7463 3187 7497
rect 3153 7395 3187 7429
rect 3153 7327 3187 7361
rect 3153 7259 3187 7293
rect 3153 7191 3187 7225
rect 3153 7123 3187 7157
rect 3153 7055 3187 7089
rect 3153 6987 3187 7021
rect 3153 6919 3187 6953
rect 3153 6851 3187 6885
rect 3153 6783 3187 6817
rect 3153 6715 3187 6749
rect 3153 6647 3187 6681
rect 3153 6579 3187 6613
rect 3153 6511 3187 6545
rect 3153 6443 3187 6477
rect 3153 6375 3187 6409
rect 3153 6307 3187 6341
rect 3153 6239 3187 6273
rect 3153 6171 3187 6205
rect 3153 6103 3187 6137
rect 3153 6035 3187 6069
rect 3153 5967 3187 6001
rect 3153 5899 3187 5933
rect 3153 5831 3187 5865
rect 3153 5763 3187 5797
rect 3153 5695 3187 5729
rect 3153 5627 3187 5661
rect 3153 5559 3187 5593
rect 3153 5491 3187 5525
rect 3153 5423 3187 5457
rect 3153 5355 3187 5389
rect 3153 5287 3187 5321
rect 3153 5219 3187 5253
rect 3153 5151 3187 5185
rect 3153 5083 3187 5117
rect 3153 5015 3187 5049
rect 3153 4947 3187 4981
rect 3153 4879 3187 4913
rect 3153 4811 3187 4845
rect 3153 4743 3187 4777
rect 3153 4675 3187 4709
rect 3153 4607 3187 4641
rect 3153 4539 3187 4573
rect 3153 4471 3187 4505
rect 3153 4403 3187 4437
rect 3153 4335 3187 4369
rect 3153 4267 3187 4301
rect 3153 4199 3187 4233
rect 3153 4131 3187 4165
rect 3153 4063 3187 4097
rect 3153 3995 3187 4029
rect 3153 3927 3187 3961
rect 3153 3859 3187 3893
rect 3153 3791 3187 3825
rect 3153 3723 3187 3757
rect 3153 3655 3187 3689
rect 3153 3587 3187 3621
rect 3153 3519 3187 3553
rect 3153 3451 3187 3485
rect 3153 3383 3187 3417
rect 3153 3315 3187 3349
rect 3153 3247 3187 3281
rect 3153 3179 3187 3213
rect 3153 3111 3187 3145
rect 3153 3043 3187 3077
rect 3153 2975 3187 3009
rect 3153 2907 3187 2941
rect 3153 2839 3187 2873
rect 3153 2771 3187 2805
rect 3153 2703 3187 2737
rect 3153 2635 3187 2669
rect 3153 2567 3187 2601
rect 3153 2499 3187 2533
rect 3153 2431 3187 2465
rect 3153 2363 3187 2397
rect 3153 2295 3187 2329
rect 3153 2227 3187 2261
rect 3153 2159 3187 2193
rect 3153 2091 3187 2125
rect 3153 2023 3187 2057
rect 3153 1955 3187 1989
rect 3153 1887 3187 1921
rect 3153 1819 3187 1853
rect 3153 1751 3187 1785
rect 3153 1683 3187 1717
rect 3153 1615 3187 1649
rect 3153 1547 3187 1581
rect 3153 1479 3187 1513
rect 3153 1411 3187 1445
rect 3153 1343 3187 1377
rect 3153 1275 3187 1309
rect 3153 1207 3187 1241
rect 3153 1139 3187 1173
rect 3153 1071 3187 1105
rect 3153 1003 3187 1037
rect 3153 935 3187 969
rect 3153 867 3187 901
rect 3153 799 3187 833
rect 3153 731 3187 765
rect 3153 663 3187 697
rect 3153 595 3187 629
rect 3153 527 3187 561
rect 3153 459 3187 493
rect 3153 391 3187 425
rect 3153 323 3187 357
rect 3153 255 3187 289
rect 3153 187 3187 221
rect 3153 119 3187 153
rect 3153 51 3187 85
rect 3153 -17 3187 17
rect 3153 -85 3187 -51
rect 3153 -153 3187 -119
rect 3153 -221 3187 -187
rect 3153 -289 3187 -255
rect 3153 -357 3187 -323
rect 3153 -425 3187 -391
rect 3153 -493 3187 -459
rect 3153 -561 3187 -527
rect 3153 -629 3187 -595
rect 3153 -697 3187 -663
rect 3153 -765 3187 -731
rect 3153 -833 3187 -799
rect 3153 -901 3187 -867
rect 3153 -969 3187 -935
rect 3153 -1037 3187 -1003
rect 3153 -1105 3187 -1071
rect 3153 -1173 3187 -1139
rect 3153 -1241 3187 -1207
rect 3153 -1309 3187 -1275
rect 3153 -1377 3187 -1343
rect 3153 -1445 3187 -1411
rect 3153 -1513 3187 -1479
rect 3153 -1581 3187 -1547
rect 3153 -1649 3187 -1615
rect 3153 -1717 3187 -1683
rect 3153 -1785 3187 -1751
rect 3153 -1853 3187 -1819
rect 3153 -1921 3187 -1887
rect 3153 -1989 3187 -1955
rect 3153 -2057 3187 -2023
rect 3153 -2125 3187 -2091
rect 3153 -2193 3187 -2159
rect 3153 -2261 3187 -2227
rect 3153 -2329 3187 -2295
rect 3153 -2397 3187 -2363
rect 3153 -2465 3187 -2431
rect 3153 -2533 3187 -2499
rect 3153 -2601 3187 -2567
rect 3153 -2669 3187 -2635
rect 3153 -2737 3187 -2703
rect 3153 -2805 3187 -2771
rect 3153 -2873 3187 -2839
rect 3153 -2941 3187 -2907
rect 3153 -3009 3187 -2975
rect 3153 -3077 3187 -3043
rect 3153 -3145 3187 -3111
rect 3153 -3213 3187 -3179
rect 3153 -3281 3187 -3247
rect 3153 -3349 3187 -3315
rect 3153 -3417 3187 -3383
rect 3153 -3485 3187 -3451
rect 3153 -3553 3187 -3519
rect 3153 -3621 3187 -3587
rect 3153 -3689 3187 -3655
rect 3153 -3757 3187 -3723
rect 3153 -3825 3187 -3791
rect 3153 -3893 3187 -3859
rect 3153 -3961 3187 -3927
rect 3153 -4029 3187 -3995
rect 3153 -4097 3187 -4063
rect 3153 -4165 3187 -4131
rect 3153 -4233 3187 -4199
rect 3153 -4301 3187 -4267
rect 3153 -4369 3187 -4335
rect 3153 -4437 3187 -4403
rect 3153 -4505 3187 -4471
rect 3153 -4573 3187 -4539
rect 3153 -4641 3187 -4607
rect 3153 -4709 3187 -4675
rect 3153 -4777 3187 -4743
rect 3153 -4845 3187 -4811
rect 3153 -4913 3187 -4879
rect 3153 -4981 3187 -4947
rect 3153 -5049 3187 -5015
rect 3153 -5117 3187 -5083
rect 3153 -5185 3187 -5151
rect 3153 -5253 3187 -5219
rect 3153 -5321 3187 -5287
rect 3153 -5389 3187 -5355
rect 3153 -5457 3187 -5423
rect 3153 -5525 3187 -5491
rect 3153 -5593 3187 -5559
rect 3153 -5661 3187 -5627
rect 3153 -5729 3187 -5695
rect 3153 -5797 3187 -5763
rect 3153 -5865 3187 -5831
rect 3153 -5933 3187 -5899
rect 3153 -6001 3187 -5967
rect 3153 -6069 3187 -6035
rect 3153 -6137 3187 -6103
rect 3153 -6205 3187 -6171
rect 3153 -6273 3187 -6239
rect 3153 -6341 3187 -6307
rect 3153 -6409 3187 -6375
rect 3153 -6477 3187 -6443
rect 3153 -6545 3187 -6511
rect 3153 -6613 3187 -6579
rect 3153 -6681 3187 -6647
rect 3153 -6749 3187 -6715
rect 3153 -6817 3187 -6783
rect 3153 -6885 3187 -6851
rect 3153 -6953 3187 -6919
rect 3153 -7021 3187 -6987
rect 3153 -7089 3187 -7055
rect 3153 -7157 3187 -7123
rect 3153 -7225 3187 -7191
rect 3153 -7293 3187 -7259
rect 3153 -7361 3187 -7327
rect 3153 -7429 3187 -7395
rect 3153 -7497 3187 -7463
rect 3153 -7565 3187 -7531
rect 3153 -7633 3187 -7599
rect 3153 -7701 3187 -7667
rect 3153 -7769 3187 -7735
rect 3153 -7837 3187 -7803
rect 3153 -7905 3187 -7871
rect 3153 -7973 3187 -7939
rect 3153 -8041 3187 -8007
rect 3153 -8109 3187 -8075
rect 3153 -8177 3187 -8143
rect 3153 -8245 3187 -8211
rect 3153 -8313 3187 -8279
rect 3153 -8381 3187 -8347
rect 3153 -8449 3187 -8415
rect 3153 -8517 3187 -8483
rect 3153 -8585 3187 -8551
rect 3153 -8653 3187 -8619
rect 3153 -8721 3187 -8687
rect 3153 -8789 3187 -8755
rect 3153 -8857 3187 -8823
rect 3153 -8925 3187 -8891
rect 3153 -8993 3187 -8959
rect 3153 -9061 3187 -9027
rect 3153 -9129 3187 -9095
rect 3153 -9197 3187 -9163
rect 3153 -9265 3187 -9231
rect 3153 -9333 3187 -9299
rect 3153 -9401 3187 -9367
rect 3153 -9469 3187 -9435
rect 3153 -9537 3187 -9503
rect 3153 -9605 3187 -9571
rect 3153 -9673 3187 -9639
rect 3153 -9741 3187 -9707
rect 3153 -9809 3187 -9775
rect 3153 -9877 3187 -9843
rect 3153 -9945 3187 -9911
rect 3153 -10013 3187 -9979
rect 3153 -10081 3187 -10047
rect 3153 -10149 3187 -10115
rect 3153 -10217 3187 -10183
rect 3153 -10285 3187 -10251
rect 3153 -10353 3187 -10319
rect 3153 -10421 3187 -10387
rect 3153 -10489 3187 -10455
rect 3153 -10557 3187 -10523
rect 3153 -10625 3187 -10591
rect 3153 -10693 3187 -10659
rect 3153 -10761 3187 -10727
rect 3153 -10829 3187 -10795
rect 3153 -10897 3187 -10863
rect 3153 -10965 3187 -10931
rect 3153 -11033 3187 -10999
rect -3077 -11162 -3043 -11128
rect -3009 -11162 -2975 -11128
rect -2941 -11162 -2907 -11128
rect -2873 -11162 -2839 -11128
rect -2805 -11162 -2771 -11128
rect -2737 -11162 -2703 -11128
rect -2669 -11162 -2635 -11128
rect -2601 -11162 -2567 -11128
rect -2533 -11162 -2499 -11128
rect -2465 -11162 -2431 -11128
rect -2397 -11162 -2363 -11128
rect -2329 -11162 -2295 -11128
rect -2261 -11162 -2227 -11128
rect -2193 -11162 -2159 -11128
rect -2125 -11162 -2091 -11128
rect -2057 -11162 -2023 -11128
rect -1989 -11162 -1955 -11128
rect -1921 -11162 -1887 -11128
rect -1853 -11162 -1819 -11128
rect -1785 -11162 -1751 -11128
rect -1717 -11162 -1683 -11128
rect -1649 -11162 -1615 -11128
rect -1581 -11162 -1547 -11128
rect -1513 -11162 -1479 -11128
rect -1445 -11162 -1411 -11128
rect -1377 -11162 -1343 -11128
rect -1309 -11162 -1275 -11128
rect -1241 -11162 -1207 -11128
rect -1173 -11162 -1139 -11128
rect -1105 -11162 -1071 -11128
rect -1037 -11162 -1003 -11128
rect -969 -11162 -935 -11128
rect -901 -11162 -867 -11128
rect -833 -11162 -799 -11128
rect -765 -11162 -731 -11128
rect -697 -11162 -663 -11128
rect -629 -11162 -595 -11128
rect -561 -11162 -527 -11128
rect -493 -11162 -459 -11128
rect -425 -11162 -391 -11128
rect -357 -11162 -323 -11128
rect -289 -11162 -255 -11128
rect -221 -11162 -187 -11128
rect -153 -11162 -119 -11128
rect -85 -11162 -51 -11128
rect -17 -11162 17 -11128
rect 51 -11162 85 -11128
rect 119 -11162 153 -11128
rect 187 -11162 221 -11128
rect 255 -11162 289 -11128
rect 323 -11162 357 -11128
rect 391 -11162 425 -11128
rect 459 -11162 493 -11128
rect 527 -11162 561 -11128
rect 595 -11162 629 -11128
rect 663 -11162 697 -11128
rect 731 -11162 765 -11128
rect 799 -11162 833 -11128
rect 867 -11162 901 -11128
rect 935 -11162 969 -11128
rect 1003 -11162 1037 -11128
rect 1071 -11162 1105 -11128
rect 1139 -11162 1173 -11128
rect 1207 -11162 1241 -11128
rect 1275 -11162 1309 -11128
rect 1343 -11162 1377 -11128
rect 1411 -11162 1445 -11128
rect 1479 -11162 1513 -11128
rect 1547 -11162 1581 -11128
rect 1615 -11162 1649 -11128
rect 1683 -11162 1717 -11128
rect 1751 -11162 1785 -11128
rect 1819 -11162 1853 -11128
rect 1887 -11162 1921 -11128
rect 1955 -11162 1989 -11128
rect 2023 -11162 2057 -11128
rect 2091 -11162 2125 -11128
rect 2159 -11162 2193 -11128
rect 2227 -11162 2261 -11128
rect 2295 -11162 2329 -11128
rect 2363 -11162 2397 -11128
rect 2431 -11162 2465 -11128
rect 2499 -11162 2533 -11128
rect 2567 -11162 2601 -11128
rect 2635 -11162 2669 -11128
rect 2703 -11162 2737 -11128
rect 2771 -11162 2805 -11128
rect 2839 -11162 2873 -11128
rect 2907 -11162 2941 -11128
rect 2975 -11162 3009 -11128
rect 3043 -11162 3077 -11128
<< xpolycontact >>
rect -3057 10600 -1911 11032
rect -3057 -11032 -1911 -10600
rect -1815 10600 -669 11032
rect -1815 -11032 -669 -10600
rect -573 10600 573 11032
rect -573 -11032 573 -10600
rect 669 10600 1815 11032
rect 669 -11032 1815 -10600
rect 1911 10600 3057 11032
rect 1911 -11032 3057 -10600
<< xpolyres >>
rect -3057 -10600 -1911 10600
rect -1815 -10600 -669 10600
rect -573 -10600 573 10600
rect 669 -10600 1815 10600
rect 1911 -10600 3057 10600
<< locali >>
rect -3187 11128 -3077 11162
rect -3043 11128 -3009 11162
rect -2975 11128 -2941 11162
rect -2907 11128 -2873 11162
rect -2839 11128 -2805 11162
rect -2771 11128 -2737 11162
rect -2703 11128 -2669 11162
rect -2635 11128 -2601 11162
rect -2567 11128 -2533 11162
rect -2499 11128 -2465 11162
rect -2431 11128 -2397 11162
rect -2363 11128 -2329 11162
rect -2295 11128 -2261 11162
rect -2227 11128 -2193 11162
rect -2159 11128 -2125 11162
rect -2091 11128 -2057 11162
rect -2023 11128 -1989 11162
rect -1955 11128 -1921 11162
rect -1887 11128 -1853 11162
rect -1819 11128 -1785 11162
rect -1751 11128 -1717 11162
rect -1683 11128 -1649 11162
rect -1615 11128 -1581 11162
rect -1547 11128 -1513 11162
rect -1479 11128 -1445 11162
rect -1411 11128 -1377 11162
rect -1343 11128 -1309 11162
rect -1275 11128 -1241 11162
rect -1207 11128 -1173 11162
rect -1139 11128 -1105 11162
rect -1071 11128 -1037 11162
rect -1003 11128 -969 11162
rect -935 11128 -901 11162
rect -867 11128 -833 11162
rect -799 11128 -765 11162
rect -731 11128 -697 11162
rect -663 11128 -629 11162
rect -595 11128 -561 11162
rect -527 11128 -493 11162
rect -459 11128 -425 11162
rect -391 11128 -357 11162
rect -323 11128 -289 11162
rect -255 11128 -221 11162
rect -187 11128 -153 11162
rect -119 11128 -85 11162
rect -51 11128 -17 11162
rect 17 11128 51 11162
rect 85 11128 119 11162
rect 153 11128 187 11162
rect 221 11128 255 11162
rect 289 11128 323 11162
rect 357 11128 391 11162
rect 425 11128 459 11162
rect 493 11128 527 11162
rect 561 11128 595 11162
rect 629 11128 663 11162
rect 697 11128 731 11162
rect 765 11128 799 11162
rect 833 11128 867 11162
rect 901 11128 935 11162
rect 969 11128 1003 11162
rect 1037 11128 1071 11162
rect 1105 11128 1139 11162
rect 1173 11128 1207 11162
rect 1241 11128 1275 11162
rect 1309 11128 1343 11162
rect 1377 11128 1411 11162
rect 1445 11128 1479 11162
rect 1513 11128 1547 11162
rect 1581 11128 1615 11162
rect 1649 11128 1683 11162
rect 1717 11128 1751 11162
rect 1785 11128 1819 11162
rect 1853 11128 1887 11162
rect 1921 11128 1955 11162
rect 1989 11128 2023 11162
rect 2057 11128 2091 11162
rect 2125 11128 2159 11162
rect 2193 11128 2227 11162
rect 2261 11128 2295 11162
rect 2329 11128 2363 11162
rect 2397 11128 2431 11162
rect 2465 11128 2499 11162
rect 2533 11128 2567 11162
rect 2601 11128 2635 11162
rect 2669 11128 2703 11162
rect 2737 11128 2771 11162
rect 2805 11128 2839 11162
rect 2873 11128 2907 11162
rect 2941 11128 2975 11162
rect 3009 11128 3043 11162
rect 3077 11128 3187 11162
rect -3187 11033 -3153 11128
rect 3153 11033 3187 11128
rect -3187 10965 -3153 10999
rect -3187 10897 -3153 10931
rect -3187 10829 -3153 10863
rect -3187 10761 -3153 10795
rect -3187 10693 -3153 10727
rect -3187 10625 -3153 10659
rect 3153 10965 3187 10999
rect 3153 10897 3187 10931
rect 3153 10829 3187 10863
rect 3153 10761 3187 10795
rect 3153 10693 3187 10727
rect 3153 10625 3187 10659
rect -3187 10557 -3153 10591
rect -3187 10489 -3153 10523
rect -3187 10421 -3153 10455
rect -3187 10353 -3153 10387
rect -3187 10285 -3153 10319
rect -3187 10217 -3153 10251
rect -3187 10149 -3153 10183
rect -3187 10081 -3153 10115
rect -3187 10013 -3153 10047
rect -3187 9945 -3153 9979
rect -3187 9877 -3153 9911
rect -3187 9809 -3153 9843
rect -3187 9741 -3153 9775
rect -3187 9673 -3153 9707
rect -3187 9605 -3153 9639
rect -3187 9537 -3153 9571
rect -3187 9469 -3153 9503
rect -3187 9401 -3153 9435
rect -3187 9333 -3153 9367
rect -3187 9265 -3153 9299
rect -3187 9197 -3153 9231
rect -3187 9129 -3153 9163
rect -3187 9061 -3153 9095
rect -3187 8993 -3153 9027
rect -3187 8925 -3153 8959
rect -3187 8857 -3153 8891
rect -3187 8789 -3153 8823
rect -3187 8721 -3153 8755
rect -3187 8653 -3153 8687
rect -3187 8585 -3153 8619
rect -3187 8517 -3153 8551
rect -3187 8449 -3153 8483
rect -3187 8381 -3153 8415
rect -3187 8313 -3153 8347
rect -3187 8245 -3153 8279
rect -3187 8177 -3153 8211
rect -3187 8109 -3153 8143
rect -3187 8041 -3153 8075
rect -3187 7973 -3153 8007
rect -3187 7905 -3153 7939
rect -3187 7837 -3153 7871
rect -3187 7769 -3153 7803
rect -3187 7701 -3153 7735
rect -3187 7633 -3153 7667
rect -3187 7565 -3153 7599
rect -3187 7497 -3153 7531
rect -3187 7429 -3153 7463
rect -3187 7361 -3153 7395
rect -3187 7293 -3153 7327
rect -3187 7225 -3153 7259
rect -3187 7157 -3153 7191
rect -3187 7089 -3153 7123
rect -3187 7021 -3153 7055
rect -3187 6953 -3153 6987
rect -3187 6885 -3153 6919
rect -3187 6817 -3153 6851
rect -3187 6749 -3153 6783
rect -3187 6681 -3153 6715
rect -3187 6613 -3153 6647
rect -3187 6545 -3153 6579
rect -3187 6477 -3153 6511
rect -3187 6409 -3153 6443
rect -3187 6341 -3153 6375
rect -3187 6273 -3153 6307
rect -3187 6205 -3153 6239
rect -3187 6137 -3153 6171
rect -3187 6069 -3153 6103
rect -3187 6001 -3153 6035
rect -3187 5933 -3153 5967
rect -3187 5865 -3153 5899
rect -3187 5797 -3153 5831
rect -3187 5729 -3153 5763
rect -3187 5661 -3153 5695
rect -3187 5593 -3153 5627
rect -3187 5525 -3153 5559
rect -3187 5457 -3153 5491
rect -3187 5389 -3153 5423
rect -3187 5321 -3153 5355
rect -3187 5253 -3153 5287
rect -3187 5185 -3153 5219
rect -3187 5117 -3153 5151
rect -3187 5049 -3153 5083
rect -3187 4981 -3153 5015
rect -3187 4913 -3153 4947
rect -3187 4845 -3153 4879
rect -3187 4777 -3153 4811
rect -3187 4709 -3153 4743
rect -3187 4641 -3153 4675
rect -3187 4573 -3153 4607
rect -3187 4505 -3153 4539
rect -3187 4437 -3153 4471
rect -3187 4369 -3153 4403
rect -3187 4301 -3153 4335
rect -3187 4233 -3153 4267
rect -3187 4165 -3153 4199
rect -3187 4097 -3153 4131
rect -3187 4029 -3153 4063
rect -3187 3961 -3153 3995
rect -3187 3893 -3153 3927
rect -3187 3825 -3153 3859
rect -3187 3757 -3153 3791
rect -3187 3689 -3153 3723
rect -3187 3621 -3153 3655
rect -3187 3553 -3153 3587
rect -3187 3485 -3153 3519
rect -3187 3417 -3153 3451
rect -3187 3349 -3153 3383
rect -3187 3281 -3153 3315
rect -3187 3213 -3153 3247
rect -3187 3145 -3153 3179
rect -3187 3077 -3153 3111
rect -3187 3009 -3153 3043
rect -3187 2941 -3153 2975
rect -3187 2873 -3153 2907
rect -3187 2805 -3153 2839
rect -3187 2737 -3153 2771
rect -3187 2669 -3153 2703
rect -3187 2601 -3153 2635
rect -3187 2533 -3153 2567
rect -3187 2465 -3153 2499
rect -3187 2397 -3153 2431
rect -3187 2329 -3153 2363
rect -3187 2261 -3153 2295
rect -3187 2193 -3153 2227
rect -3187 2125 -3153 2159
rect -3187 2057 -3153 2091
rect -3187 1989 -3153 2023
rect -3187 1921 -3153 1955
rect -3187 1853 -3153 1887
rect -3187 1785 -3153 1819
rect -3187 1717 -3153 1751
rect -3187 1649 -3153 1683
rect -3187 1581 -3153 1615
rect -3187 1513 -3153 1547
rect -3187 1445 -3153 1479
rect -3187 1377 -3153 1411
rect -3187 1309 -3153 1343
rect -3187 1241 -3153 1275
rect -3187 1173 -3153 1207
rect -3187 1105 -3153 1139
rect -3187 1037 -3153 1071
rect -3187 969 -3153 1003
rect -3187 901 -3153 935
rect -3187 833 -3153 867
rect -3187 765 -3153 799
rect -3187 697 -3153 731
rect -3187 629 -3153 663
rect -3187 561 -3153 595
rect -3187 493 -3153 527
rect -3187 425 -3153 459
rect -3187 357 -3153 391
rect -3187 289 -3153 323
rect -3187 221 -3153 255
rect -3187 153 -3153 187
rect -3187 85 -3153 119
rect -3187 17 -3153 51
rect -3187 -51 -3153 -17
rect -3187 -119 -3153 -85
rect -3187 -187 -3153 -153
rect -3187 -255 -3153 -221
rect -3187 -323 -3153 -289
rect -3187 -391 -3153 -357
rect -3187 -459 -3153 -425
rect -3187 -527 -3153 -493
rect -3187 -595 -3153 -561
rect -3187 -663 -3153 -629
rect -3187 -731 -3153 -697
rect -3187 -799 -3153 -765
rect -3187 -867 -3153 -833
rect -3187 -935 -3153 -901
rect -3187 -1003 -3153 -969
rect -3187 -1071 -3153 -1037
rect -3187 -1139 -3153 -1105
rect -3187 -1207 -3153 -1173
rect -3187 -1275 -3153 -1241
rect -3187 -1343 -3153 -1309
rect -3187 -1411 -3153 -1377
rect -3187 -1479 -3153 -1445
rect -3187 -1547 -3153 -1513
rect -3187 -1615 -3153 -1581
rect -3187 -1683 -3153 -1649
rect -3187 -1751 -3153 -1717
rect -3187 -1819 -3153 -1785
rect -3187 -1887 -3153 -1853
rect -3187 -1955 -3153 -1921
rect -3187 -2023 -3153 -1989
rect -3187 -2091 -3153 -2057
rect -3187 -2159 -3153 -2125
rect -3187 -2227 -3153 -2193
rect -3187 -2295 -3153 -2261
rect -3187 -2363 -3153 -2329
rect -3187 -2431 -3153 -2397
rect -3187 -2499 -3153 -2465
rect -3187 -2567 -3153 -2533
rect -3187 -2635 -3153 -2601
rect -3187 -2703 -3153 -2669
rect -3187 -2771 -3153 -2737
rect -3187 -2839 -3153 -2805
rect -3187 -2907 -3153 -2873
rect -3187 -2975 -3153 -2941
rect -3187 -3043 -3153 -3009
rect -3187 -3111 -3153 -3077
rect -3187 -3179 -3153 -3145
rect -3187 -3247 -3153 -3213
rect -3187 -3315 -3153 -3281
rect -3187 -3383 -3153 -3349
rect -3187 -3451 -3153 -3417
rect -3187 -3519 -3153 -3485
rect -3187 -3587 -3153 -3553
rect -3187 -3655 -3153 -3621
rect -3187 -3723 -3153 -3689
rect -3187 -3791 -3153 -3757
rect -3187 -3859 -3153 -3825
rect -3187 -3927 -3153 -3893
rect -3187 -3995 -3153 -3961
rect -3187 -4063 -3153 -4029
rect -3187 -4131 -3153 -4097
rect -3187 -4199 -3153 -4165
rect -3187 -4267 -3153 -4233
rect -3187 -4335 -3153 -4301
rect -3187 -4403 -3153 -4369
rect -3187 -4471 -3153 -4437
rect -3187 -4539 -3153 -4505
rect -3187 -4607 -3153 -4573
rect -3187 -4675 -3153 -4641
rect -3187 -4743 -3153 -4709
rect -3187 -4811 -3153 -4777
rect -3187 -4879 -3153 -4845
rect -3187 -4947 -3153 -4913
rect -3187 -5015 -3153 -4981
rect -3187 -5083 -3153 -5049
rect -3187 -5151 -3153 -5117
rect -3187 -5219 -3153 -5185
rect -3187 -5287 -3153 -5253
rect -3187 -5355 -3153 -5321
rect -3187 -5423 -3153 -5389
rect -3187 -5491 -3153 -5457
rect -3187 -5559 -3153 -5525
rect -3187 -5627 -3153 -5593
rect -3187 -5695 -3153 -5661
rect -3187 -5763 -3153 -5729
rect -3187 -5831 -3153 -5797
rect -3187 -5899 -3153 -5865
rect -3187 -5967 -3153 -5933
rect -3187 -6035 -3153 -6001
rect -3187 -6103 -3153 -6069
rect -3187 -6171 -3153 -6137
rect -3187 -6239 -3153 -6205
rect -3187 -6307 -3153 -6273
rect -3187 -6375 -3153 -6341
rect -3187 -6443 -3153 -6409
rect -3187 -6511 -3153 -6477
rect -3187 -6579 -3153 -6545
rect -3187 -6647 -3153 -6613
rect -3187 -6715 -3153 -6681
rect -3187 -6783 -3153 -6749
rect -3187 -6851 -3153 -6817
rect -3187 -6919 -3153 -6885
rect -3187 -6987 -3153 -6953
rect -3187 -7055 -3153 -7021
rect -3187 -7123 -3153 -7089
rect -3187 -7191 -3153 -7157
rect -3187 -7259 -3153 -7225
rect -3187 -7327 -3153 -7293
rect -3187 -7395 -3153 -7361
rect -3187 -7463 -3153 -7429
rect -3187 -7531 -3153 -7497
rect -3187 -7599 -3153 -7565
rect -3187 -7667 -3153 -7633
rect -3187 -7735 -3153 -7701
rect -3187 -7803 -3153 -7769
rect -3187 -7871 -3153 -7837
rect -3187 -7939 -3153 -7905
rect -3187 -8007 -3153 -7973
rect -3187 -8075 -3153 -8041
rect -3187 -8143 -3153 -8109
rect -3187 -8211 -3153 -8177
rect -3187 -8279 -3153 -8245
rect -3187 -8347 -3153 -8313
rect -3187 -8415 -3153 -8381
rect -3187 -8483 -3153 -8449
rect -3187 -8551 -3153 -8517
rect -3187 -8619 -3153 -8585
rect -3187 -8687 -3153 -8653
rect -3187 -8755 -3153 -8721
rect -3187 -8823 -3153 -8789
rect -3187 -8891 -3153 -8857
rect -3187 -8959 -3153 -8925
rect -3187 -9027 -3153 -8993
rect -3187 -9095 -3153 -9061
rect -3187 -9163 -3153 -9129
rect -3187 -9231 -3153 -9197
rect -3187 -9299 -3153 -9265
rect -3187 -9367 -3153 -9333
rect -3187 -9435 -3153 -9401
rect -3187 -9503 -3153 -9469
rect -3187 -9571 -3153 -9537
rect -3187 -9639 -3153 -9605
rect -3187 -9707 -3153 -9673
rect -3187 -9775 -3153 -9741
rect -3187 -9843 -3153 -9809
rect -3187 -9911 -3153 -9877
rect -3187 -9979 -3153 -9945
rect -3187 -10047 -3153 -10013
rect -3187 -10115 -3153 -10081
rect -3187 -10183 -3153 -10149
rect -3187 -10251 -3153 -10217
rect -3187 -10319 -3153 -10285
rect -3187 -10387 -3153 -10353
rect -3187 -10455 -3153 -10421
rect -3187 -10523 -3153 -10489
rect -3187 -10591 -3153 -10557
rect 3153 10557 3187 10591
rect 3153 10489 3187 10523
rect 3153 10421 3187 10455
rect 3153 10353 3187 10387
rect 3153 10285 3187 10319
rect 3153 10217 3187 10251
rect 3153 10149 3187 10183
rect 3153 10081 3187 10115
rect 3153 10013 3187 10047
rect 3153 9945 3187 9979
rect 3153 9877 3187 9911
rect 3153 9809 3187 9843
rect 3153 9741 3187 9775
rect 3153 9673 3187 9707
rect 3153 9605 3187 9639
rect 3153 9537 3187 9571
rect 3153 9469 3187 9503
rect 3153 9401 3187 9435
rect 3153 9333 3187 9367
rect 3153 9265 3187 9299
rect 3153 9197 3187 9231
rect 3153 9129 3187 9163
rect 3153 9061 3187 9095
rect 3153 8993 3187 9027
rect 3153 8925 3187 8959
rect 3153 8857 3187 8891
rect 3153 8789 3187 8823
rect 3153 8721 3187 8755
rect 3153 8653 3187 8687
rect 3153 8585 3187 8619
rect 3153 8517 3187 8551
rect 3153 8449 3187 8483
rect 3153 8381 3187 8415
rect 3153 8313 3187 8347
rect 3153 8245 3187 8279
rect 3153 8177 3187 8211
rect 3153 8109 3187 8143
rect 3153 8041 3187 8075
rect 3153 7973 3187 8007
rect 3153 7905 3187 7939
rect 3153 7837 3187 7871
rect 3153 7769 3187 7803
rect 3153 7701 3187 7735
rect 3153 7633 3187 7667
rect 3153 7565 3187 7599
rect 3153 7497 3187 7531
rect 3153 7429 3187 7463
rect 3153 7361 3187 7395
rect 3153 7293 3187 7327
rect 3153 7225 3187 7259
rect 3153 7157 3187 7191
rect 3153 7089 3187 7123
rect 3153 7021 3187 7055
rect 3153 6953 3187 6987
rect 3153 6885 3187 6919
rect 3153 6817 3187 6851
rect 3153 6749 3187 6783
rect 3153 6681 3187 6715
rect 3153 6613 3187 6647
rect 3153 6545 3187 6579
rect 3153 6477 3187 6511
rect 3153 6409 3187 6443
rect 3153 6341 3187 6375
rect 3153 6273 3187 6307
rect 3153 6205 3187 6239
rect 3153 6137 3187 6171
rect 3153 6069 3187 6103
rect 3153 6001 3187 6035
rect 3153 5933 3187 5967
rect 3153 5865 3187 5899
rect 3153 5797 3187 5831
rect 3153 5729 3187 5763
rect 3153 5661 3187 5695
rect 3153 5593 3187 5627
rect 3153 5525 3187 5559
rect 3153 5457 3187 5491
rect 3153 5389 3187 5423
rect 3153 5321 3187 5355
rect 3153 5253 3187 5287
rect 3153 5185 3187 5219
rect 3153 5117 3187 5151
rect 3153 5049 3187 5083
rect 3153 4981 3187 5015
rect 3153 4913 3187 4947
rect 3153 4845 3187 4879
rect 3153 4777 3187 4811
rect 3153 4709 3187 4743
rect 3153 4641 3187 4675
rect 3153 4573 3187 4607
rect 3153 4505 3187 4539
rect 3153 4437 3187 4471
rect 3153 4369 3187 4403
rect 3153 4301 3187 4335
rect 3153 4233 3187 4267
rect 3153 4165 3187 4199
rect 3153 4097 3187 4131
rect 3153 4029 3187 4063
rect 3153 3961 3187 3995
rect 3153 3893 3187 3927
rect 3153 3825 3187 3859
rect 3153 3757 3187 3791
rect 3153 3689 3187 3723
rect 3153 3621 3187 3655
rect 3153 3553 3187 3587
rect 3153 3485 3187 3519
rect 3153 3417 3187 3451
rect 3153 3349 3187 3383
rect 3153 3281 3187 3315
rect 3153 3213 3187 3247
rect 3153 3145 3187 3179
rect 3153 3077 3187 3111
rect 3153 3009 3187 3043
rect 3153 2941 3187 2975
rect 3153 2873 3187 2907
rect 3153 2805 3187 2839
rect 3153 2737 3187 2771
rect 3153 2669 3187 2703
rect 3153 2601 3187 2635
rect 3153 2533 3187 2567
rect 3153 2465 3187 2499
rect 3153 2397 3187 2431
rect 3153 2329 3187 2363
rect 3153 2261 3187 2295
rect 3153 2193 3187 2227
rect 3153 2125 3187 2159
rect 3153 2057 3187 2091
rect 3153 1989 3187 2023
rect 3153 1921 3187 1955
rect 3153 1853 3187 1887
rect 3153 1785 3187 1819
rect 3153 1717 3187 1751
rect 3153 1649 3187 1683
rect 3153 1581 3187 1615
rect 3153 1513 3187 1547
rect 3153 1445 3187 1479
rect 3153 1377 3187 1411
rect 3153 1309 3187 1343
rect 3153 1241 3187 1275
rect 3153 1173 3187 1207
rect 3153 1105 3187 1139
rect 3153 1037 3187 1071
rect 3153 969 3187 1003
rect 3153 901 3187 935
rect 3153 833 3187 867
rect 3153 765 3187 799
rect 3153 697 3187 731
rect 3153 629 3187 663
rect 3153 561 3187 595
rect 3153 493 3187 527
rect 3153 425 3187 459
rect 3153 357 3187 391
rect 3153 289 3187 323
rect 3153 221 3187 255
rect 3153 153 3187 187
rect 3153 85 3187 119
rect 3153 17 3187 51
rect 3153 -51 3187 -17
rect 3153 -119 3187 -85
rect 3153 -187 3187 -153
rect 3153 -255 3187 -221
rect 3153 -323 3187 -289
rect 3153 -391 3187 -357
rect 3153 -459 3187 -425
rect 3153 -527 3187 -493
rect 3153 -595 3187 -561
rect 3153 -663 3187 -629
rect 3153 -731 3187 -697
rect 3153 -799 3187 -765
rect 3153 -867 3187 -833
rect 3153 -935 3187 -901
rect 3153 -1003 3187 -969
rect 3153 -1071 3187 -1037
rect 3153 -1139 3187 -1105
rect 3153 -1207 3187 -1173
rect 3153 -1275 3187 -1241
rect 3153 -1343 3187 -1309
rect 3153 -1411 3187 -1377
rect 3153 -1479 3187 -1445
rect 3153 -1547 3187 -1513
rect 3153 -1615 3187 -1581
rect 3153 -1683 3187 -1649
rect 3153 -1751 3187 -1717
rect 3153 -1819 3187 -1785
rect 3153 -1887 3187 -1853
rect 3153 -1955 3187 -1921
rect 3153 -2023 3187 -1989
rect 3153 -2091 3187 -2057
rect 3153 -2159 3187 -2125
rect 3153 -2227 3187 -2193
rect 3153 -2295 3187 -2261
rect 3153 -2363 3187 -2329
rect 3153 -2431 3187 -2397
rect 3153 -2499 3187 -2465
rect 3153 -2567 3187 -2533
rect 3153 -2635 3187 -2601
rect 3153 -2703 3187 -2669
rect 3153 -2771 3187 -2737
rect 3153 -2839 3187 -2805
rect 3153 -2907 3187 -2873
rect 3153 -2975 3187 -2941
rect 3153 -3043 3187 -3009
rect 3153 -3111 3187 -3077
rect 3153 -3179 3187 -3145
rect 3153 -3247 3187 -3213
rect 3153 -3315 3187 -3281
rect 3153 -3383 3187 -3349
rect 3153 -3451 3187 -3417
rect 3153 -3519 3187 -3485
rect 3153 -3587 3187 -3553
rect 3153 -3655 3187 -3621
rect 3153 -3723 3187 -3689
rect 3153 -3791 3187 -3757
rect 3153 -3859 3187 -3825
rect 3153 -3927 3187 -3893
rect 3153 -3995 3187 -3961
rect 3153 -4063 3187 -4029
rect 3153 -4131 3187 -4097
rect 3153 -4199 3187 -4165
rect 3153 -4267 3187 -4233
rect 3153 -4335 3187 -4301
rect 3153 -4403 3187 -4369
rect 3153 -4471 3187 -4437
rect 3153 -4539 3187 -4505
rect 3153 -4607 3187 -4573
rect 3153 -4675 3187 -4641
rect 3153 -4743 3187 -4709
rect 3153 -4811 3187 -4777
rect 3153 -4879 3187 -4845
rect 3153 -4947 3187 -4913
rect 3153 -5015 3187 -4981
rect 3153 -5083 3187 -5049
rect 3153 -5151 3187 -5117
rect 3153 -5219 3187 -5185
rect 3153 -5287 3187 -5253
rect 3153 -5355 3187 -5321
rect 3153 -5423 3187 -5389
rect 3153 -5491 3187 -5457
rect 3153 -5559 3187 -5525
rect 3153 -5627 3187 -5593
rect 3153 -5695 3187 -5661
rect 3153 -5763 3187 -5729
rect 3153 -5831 3187 -5797
rect 3153 -5899 3187 -5865
rect 3153 -5967 3187 -5933
rect 3153 -6035 3187 -6001
rect 3153 -6103 3187 -6069
rect 3153 -6171 3187 -6137
rect 3153 -6239 3187 -6205
rect 3153 -6307 3187 -6273
rect 3153 -6375 3187 -6341
rect 3153 -6443 3187 -6409
rect 3153 -6511 3187 -6477
rect 3153 -6579 3187 -6545
rect 3153 -6647 3187 -6613
rect 3153 -6715 3187 -6681
rect 3153 -6783 3187 -6749
rect 3153 -6851 3187 -6817
rect 3153 -6919 3187 -6885
rect 3153 -6987 3187 -6953
rect 3153 -7055 3187 -7021
rect 3153 -7123 3187 -7089
rect 3153 -7191 3187 -7157
rect 3153 -7259 3187 -7225
rect 3153 -7327 3187 -7293
rect 3153 -7395 3187 -7361
rect 3153 -7463 3187 -7429
rect 3153 -7531 3187 -7497
rect 3153 -7599 3187 -7565
rect 3153 -7667 3187 -7633
rect 3153 -7735 3187 -7701
rect 3153 -7803 3187 -7769
rect 3153 -7871 3187 -7837
rect 3153 -7939 3187 -7905
rect 3153 -8007 3187 -7973
rect 3153 -8075 3187 -8041
rect 3153 -8143 3187 -8109
rect 3153 -8211 3187 -8177
rect 3153 -8279 3187 -8245
rect 3153 -8347 3187 -8313
rect 3153 -8415 3187 -8381
rect 3153 -8483 3187 -8449
rect 3153 -8551 3187 -8517
rect 3153 -8619 3187 -8585
rect 3153 -8687 3187 -8653
rect 3153 -8755 3187 -8721
rect 3153 -8823 3187 -8789
rect 3153 -8891 3187 -8857
rect 3153 -8959 3187 -8925
rect 3153 -9027 3187 -8993
rect 3153 -9095 3187 -9061
rect 3153 -9163 3187 -9129
rect 3153 -9231 3187 -9197
rect 3153 -9299 3187 -9265
rect 3153 -9367 3187 -9333
rect 3153 -9435 3187 -9401
rect 3153 -9503 3187 -9469
rect 3153 -9571 3187 -9537
rect 3153 -9639 3187 -9605
rect 3153 -9707 3187 -9673
rect 3153 -9775 3187 -9741
rect 3153 -9843 3187 -9809
rect 3153 -9911 3187 -9877
rect 3153 -9979 3187 -9945
rect 3153 -10047 3187 -10013
rect 3153 -10115 3187 -10081
rect 3153 -10183 3187 -10149
rect 3153 -10251 3187 -10217
rect 3153 -10319 3187 -10285
rect 3153 -10387 3187 -10353
rect 3153 -10455 3187 -10421
rect 3153 -10523 3187 -10489
rect 3153 -10591 3187 -10557
rect -3187 -10659 -3153 -10625
rect -3187 -10727 -3153 -10693
rect -3187 -10795 -3153 -10761
rect -3187 -10863 -3153 -10829
rect -3187 -10931 -3153 -10897
rect -3187 -10999 -3153 -10965
rect 3153 -10659 3187 -10625
rect 3153 -10727 3187 -10693
rect 3153 -10795 3187 -10761
rect 3153 -10863 3187 -10829
rect 3153 -10931 3187 -10897
rect 3153 -10999 3187 -10965
rect -3187 -11128 -3153 -11033
rect 3153 -11128 3187 -11033
rect -3187 -11162 -3077 -11128
rect -3043 -11162 -3009 -11128
rect -2975 -11162 -2941 -11128
rect -2907 -11162 -2873 -11128
rect -2839 -11162 -2805 -11128
rect -2771 -11162 -2737 -11128
rect -2703 -11162 -2669 -11128
rect -2635 -11162 -2601 -11128
rect -2567 -11162 -2533 -11128
rect -2499 -11162 -2465 -11128
rect -2431 -11162 -2397 -11128
rect -2363 -11162 -2329 -11128
rect -2295 -11162 -2261 -11128
rect -2227 -11162 -2193 -11128
rect -2159 -11162 -2125 -11128
rect -2091 -11162 -2057 -11128
rect -2023 -11162 -1989 -11128
rect -1955 -11162 -1921 -11128
rect -1887 -11162 -1853 -11128
rect -1819 -11162 -1785 -11128
rect -1751 -11162 -1717 -11128
rect -1683 -11162 -1649 -11128
rect -1615 -11162 -1581 -11128
rect -1547 -11162 -1513 -11128
rect -1479 -11162 -1445 -11128
rect -1411 -11162 -1377 -11128
rect -1343 -11162 -1309 -11128
rect -1275 -11162 -1241 -11128
rect -1207 -11162 -1173 -11128
rect -1139 -11162 -1105 -11128
rect -1071 -11162 -1037 -11128
rect -1003 -11162 -969 -11128
rect -935 -11162 -901 -11128
rect -867 -11162 -833 -11128
rect -799 -11162 -765 -11128
rect -731 -11162 -697 -11128
rect -663 -11162 -629 -11128
rect -595 -11162 -561 -11128
rect -527 -11162 -493 -11128
rect -459 -11162 -425 -11128
rect -391 -11162 -357 -11128
rect -323 -11162 -289 -11128
rect -255 -11162 -221 -11128
rect -187 -11162 -153 -11128
rect -119 -11162 -85 -11128
rect -51 -11162 -17 -11128
rect 17 -11162 51 -11128
rect 85 -11162 119 -11128
rect 153 -11162 187 -11128
rect 221 -11162 255 -11128
rect 289 -11162 323 -11128
rect 357 -11162 391 -11128
rect 425 -11162 459 -11128
rect 493 -11162 527 -11128
rect 561 -11162 595 -11128
rect 629 -11162 663 -11128
rect 697 -11162 731 -11128
rect 765 -11162 799 -11128
rect 833 -11162 867 -11128
rect 901 -11162 935 -11128
rect 969 -11162 1003 -11128
rect 1037 -11162 1071 -11128
rect 1105 -11162 1139 -11128
rect 1173 -11162 1207 -11128
rect 1241 -11162 1275 -11128
rect 1309 -11162 1343 -11128
rect 1377 -11162 1411 -11128
rect 1445 -11162 1479 -11128
rect 1513 -11162 1547 -11128
rect 1581 -11162 1615 -11128
rect 1649 -11162 1683 -11128
rect 1717 -11162 1751 -11128
rect 1785 -11162 1819 -11128
rect 1853 -11162 1887 -11128
rect 1921 -11162 1955 -11128
rect 1989 -11162 2023 -11128
rect 2057 -11162 2091 -11128
rect 2125 -11162 2159 -11128
rect 2193 -11162 2227 -11128
rect 2261 -11162 2295 -11128
rect 2329 -11162 2363 -11128
rect 2397 -11162 2431 -11128
rect 2465 -11162 2499 -11128
rect 2533 -11162 2567 -11128
rect 2601 -11162 2635 -11128
rect 2669 -11162 2703 -11128
rect 2737 -11162 2771 -11128
rect 2805 -11162 2839 -11128
rect 2873 -11162 2907 -11128
rect 2941 -11162 2975 -11128
rect 3009 -11162 3043 -11128
rect 3077 -11162 3187 -11128
<< viali >>
rect -3041 10618 -1927 11012
rect -1799 10618 -685 11012
rect -557 10618 557 11012
rect 685 10618 1799 11012
rect 1927 10618 3041 11012
rect -3041 -11013 -1927 -10619
rect -1799 -11013 -685 -10619
rect -557 -11013 557 -10619
rect 685 -11013 1799 -10619
rect 1927 -11013 3041 -10619
<< metal1 >>
rect -3053 11012 -1915 11020
rect -3053 10618 -3041 11012
rect -1927 10618 -1915 11012
rect -3053 10611 -1915 10618
rect -1811 11012 -673 11020
rect -1811 10618 -1799 11012
rect -685 10618 -673 11012
rect -1811 10611 -673 10618
rect -569 11012 569 11020
rect -569 10618 -557 11012
rect 557 10618 569 11012
rect -569 10611 569 10618
rect 673 11012 1811 11020
rect 673 10618 685 11012
rect 1799 10618 1811 11012
rect 673 10611 1811 10618
rect 1915 11012 3053 11020
rect 1915 10618 1927 11012
rect 3041 10618 3053 11012
rect 1915 10611 3053 10618
rect -3053 -10619 -1915 -10611
rect -3053 -11013 -3041 -10619
rect -1927 -11013 -1915 -10619
rect -3053 -11020 -1915 -11013
rect -1811 -10619 -673 -10611
rect -1811 -11013 -1799 -10619
rect -685 -11013 -673 -10619
rect -1811 -11020 -673 -11013
rect -569 -10619 569 -10611
rect -569 -11013 -557 -10619
rect 557 -11013 569 -10619
rect -569 -11020 569 -11013
rect 673 -10619 1811 -10611
rect 673 -11013 685 -10619
rect 1799 -11013 1811 -10619
rect 673 -11020 1811 -11013
rect 1915 -10619 3053 -10611
rect 1915 -11013 1927 -10619
rect 3041 -11013 3053 -10619
rect 1915 -11020 3053 -11013
<< properties >>
string FIXED_BBOX -3170 -11145 3170 11145
<< end >>
