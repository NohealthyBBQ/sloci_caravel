magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 244 5462 278 5542
rect 876 5462 910 5542
rect 1508 5462 1542 5542
rect 2140 5462 2174 5542
rect 2400 5453 2440 5470
rect 2400 5419 2403 5453
rect 2437 5419 2440 5453
rect 2400 5381 2440 5419
rect 2400 5347 2403 5381
rect 2437 5347 2440 5381
rect 2400 5330 2440 5347
rect 2400 4093 2440 4110
rect 2400 4059 2403 4093
rect 2437 4059 2440 4093
rect 2400 4021 2440 4059
rect 2400 3987 2403 4021
rect 2437 3987 2440 4021
rect 2400 3970 2440 3987
rect 2400 2723 2440 2740
rect 2400 2689 2403 2723
rect 2437 2689 2440 2723
rect 2400 2651 2440 2689
rect 2400 2617 2403 2651
rect 2437 2617 2440 2651
rect 2400 2600 2440 2617
rect 2400 1363 2440 1380
rect 2400 1329 2403 1363
rect 2437 1329 2440 1363
rect 2400 1291 2440 1329
rect 2400 1257 2403 1291
rect 2437 1257 2440 1291
rect 2400 1240 2440 1257
<< viali >>
rect 2403 5419 2437 5453
rect 2403 5347 2437 5381
rect 2403 4059 2437 4093
rect 2403 3987 2437 4021
rect 2403 2689 2437 2723
rect 2403 2617 2437 2651
rect 2403 1329 2437 1363
rect 2403 1257 2437 1291
<< metal1 >>
rect 212 5460 312 5462
rect 212 5408 236 5460
rect 288 5408 312 5460
rect 212 5396 312 5408
rect 212 5344 236 5396
rect 288 5344 312 5396
rect 212 5342 312 5344
rect 396 5449 442 5465
rect 396 4380 402 5449
rect 436 4380 442 5449
rect 528 5460 628 5462
rect 528 5408 552 5460
rect 604 5408 628 5460
rect 528 5396 628 5408
rect 528 5344 552 5396
rect 604 5344 628 5396
rect 528 5342 628 5344
rect 712 5449 758 5461
rect 52 4378 152 4380
rect 52 4326 76 4378
rect 128 4326 152 4378
rect 52 4314 152 4326
rect 52 4262 76 4314
rect 128 4262 152 4314
rect 52 4260 152 4262
rect 368 4378 468 4380
rect 368 4326 392 4378
rect 444 4326 468 4378
rect 368 4314 468 4326
rect 368 4262 392 4314
rect 444 4262 468 4314
rect 368 4260 468 4262
rect 554 4273 560 5342
rect 594 4277 600 5342
rect 712 4380 718 5449
rect 752 4380 758 5449
rect 844 5460 944 5462
rect 844 5408 868 5460
rect 920 5408 944 5460
rect 844 5396 944 5408
rect 844 5344 868 5396
rect 920 5344 944 5396
rect 844 5342 944 5344
rect 1028 5449 1074 5461
rect 568 4273 600 4277
rect 554 4261 600 4273
rect 684 4378 784 4380
rect 684 4326 708 4378
rect 760 4326 784 4378
rect 684 4314 784 4326
rect 684 4262 708 4314
rect 760 4262 784 4314
rect 684 4260 784 4262
rect 870 4273 876 5342
rect 910 4273 916 5342
rect 1028 4380 1034 5449
rect 1068 4380 1074 5449
rect 1160 5460 1260 5462
rect 1160 5408 1184 5460
rect 1236 5408 1260 5460
rect 1160 5396 1260 5408
rect 1160 5344 1184 5396
rect 1236 5344 1260 5396
rect 1160 5342 1260 5344
rect 1344 5449 1390 5465
rect 870 4261 916 4273
rect 1000 4378 1100 4380
rect 1000 4326 1024 4378
rect 1076 4326 1100 4378
rect 1000 4314 1100 4326
rect 1000 4262 1024 4314
rect 1076 4262 1100 4314
rect 1000 4260 1100 4262
rect 1186 4273 1192 5342
rect 1226 4273 1232 5342
rect 1344 4380 1350 5449
rect 1384 4380 1390 5449
rect 1476 5460 1576 5462
rect 1476 5408 1500 5460
rect 1552 5408 1576 5460
rect 1476 5396 1576 5408
rect 1476 5344 1500 5396
rect 1552 5344 1576 5396
rect 1476 5342 1576 5344
rect 1660 5449 1706 5461
rect 1186 4261 1232 4273
rect 1316 4378 1416 4380
rect 1316 4326 1340 4378
rect 1392 4326 1416 4378
rect 1316 4314 1416 4326
rect 1316 4262 1340 4314
rect 1392 4262 1416 4314
rect 1316 4260 1416 4262
rect 1502 4273 1508 5342
rect 1542 4277 1548 5342
rect 1660 4380 1666 5449
rect 1700 4380 1706 5449
rect 1792 5460 1892 5462
rect 1792 5408 1816 5460
rect 1868 5408 1892 5460
rect 1792 5396 1892 5408
rect 1792 5344 1816 5396
rect 1868 5344 1892 5396
rect 1792 5342 1892 5344
rect 1976 5449 2022 5461
rect 1516 4273 1548 4277
rect 1502 4261 1548 4273
rect 1632 4378 1732 4380
rect 1632 4326 1656 4378
rect 1708 4326 1732 4378
rect 1632 4314 1732 4326
rect 1632 4262 1656 4314
rect 1708 4262 1732 4314
rect 1632 4260 1732 4262
rect 1818 4273 1824 5342
rect 1858 4273 1864 5342
rect 1976 4380 1982 5449
rect 2016 4380 2022 5449
rect 2108 5460 2208 5462
rect 2108 5408 2132 5460
rect 2184 5408 2208 5460
rect 2108 5396 2208 5408
rect 2108 5344 2132 5396
rect 2184 5344 2208 5396
rect 2108 5342 2208 5344
rect 2292 5449 2338 5465
rect 2394 5460 2446 5482
rect 1818 4261 1864 4273
rect 1948 4378 2048 4380
rect 1948 4326 1972 4378
rect 2024 4326 2048 4378
rect 1948 4314 2048 4326
rect 1948 4262 1972 4314
rect 2024 4262 2048 4314
rect 1948 4260 2048 4262
rect 2134 4273 2140 5342
rect 2174 4273 2180 5342
rect 2292 4380 2298 5449
rect 2332 4380 2338 5449
rect 2370 5458 2450 5460
rect 2370 5406 2384 5458
rect 2436 5453 2450 5458
rect 2437 5419 2450 5453
rect 2436 5406 2450 5419
rect 2370 5394 2450 5406
rect 2370 5342 2384 5394
rect 2436 5381 2450 5394
rect 2437 5347 2450 5381
rect 2436 5342 2450 5347
rect 2370 5340 2450 5342
rect 2394 5318 2446 5340
rect 2134 4261 2180 4273
rect 2264 4378 2364 4380
rect 2264 4326 2288 4378
rect 2340 4326 2364 4378
rect 2264 4314 2364 4326
rect 2264 4262 2288 4314
rect 2340 4262 2364 4314
rect 2264 4260 2364 4262
rect -140 4214 -70 4220
rect -140 4180 142 4214
rect -140 2850 -70 4180
rect 147 4174 2293 4220
rect 80 4085 126 4097
rect 80 3016 86 4085
rect 120 3016 126 4085
rect 212 4096 312 4098
rect 212 4044 236 4096
rect 288 4044 312 4096
rect 212 4032 312 4044
rect 212 3980 236 4032
rect 288 3980 312 4032
rect 212 3978 312 3980
rect 396 4085 442 4101
rect 52 3014 152 3016
rect 52 2962 76 3014
rect 128 2962 152 3014
rect 52 2950 152 2962
rect 52 2898 76 2950
rect 128 2898 152 2950
rect 52 2896 152 2898
rect 238 2909 244 3978
rect 278 2909 284 3978
rect 396 3016 402 4085
rect 436 3016 442 4085
rect 528 4096 628 4098
rect 528 4044 552 4096
rect 604 4044 628 4096
rect 528 4032 628 4044
rect 528 3980 552 4032
rect 604 3980 628 4032
rect 528 3978 628 3980
rect 712 4085 758 4097
rect 238 2897 284 2909
rect 368 3014 468 3016
rect 368 2962 392 3014
rect 444 2962 468 3014
rect 368 2950 468 2962
rect 368 2898 392 2950
rect 444 2898 468 2950
rect 368 2896 468 2898
rect 554 2909 560 3978
rect 594 2913 600 3978
rect 712 3016 718 4085
rect 752 3016 758 4085
rect 844 4096 944 4098
rect 844 4044 868 4096
rect 920 4044 944 4096
rect 844 4032 944 4044
rect 844 3980 868 4032
rect 920 3980 944 4032
rect 844 3978 944 3980
rect 1028 4085 1074 4097
rect 568 2909 600 2913
rect 554 2897 600 2909
rect 684 3014 784 3016
rect 684 2962 708 3014
rect 760 2962 784 3014
rect 684 2950 784 2962
rect 684 2898 708 2950
rect 760 2898 784 2950
rect 684 2896 784 2898
rect 870 2909 876 3978
rect 910 2909 916 3978
rect 1028 3016 1034 4085
rect 1068 3016 1074 4085
rect 1160 4096 1260 4098
rect 1160 4044 1184 4096
rect 1236 4044 1260 4096
rect 1160 4032 1260 4044
rect 1160 3980 1184 4032
rect 1236 3980 1260 4032
rect 1160 3978 1260 3980
rect 1344 4085 1390 4101
rect 870 2897 916 2909
rect 1000 3014 1100 3016
rect 1000 2962 1024 3014
rect 1076 2962 1100 3014
rect 1000 2950 1100 2962
rect 1000 2898 1024 2950
rect 1076 2898 1100 2950
rect 1000 2896 1100 2898
rect 1186 2909 1192 3978
rect 1226 2909 1232 3978
rect 1344 3016 1350 4085
rect 1384 3016 1390 4085
rect 1476 4096 1576 4098
rect 1476 4044 1500 4096
rect 1552 4044 1576 4096
rect 1476 4032 1576 4044
rect 1476 3980 1500 4032
rect 1552 3980 1576 4032
rect 1476 3978 1576 3980
rect 1660 4085 1706 4097
rect 1186 2897 1232 2909
rect 1316 3014 1416 3016
rect 1316 2962 1340 3014
rect 1392 2962 1416 3014
rect 1316 2950 1416 2962
rect 1316 2898 1340 2950
rect 1392 2898 1416 2950
rect 1316 2896 1416 2898
rect 1502 2909 1508 3978
rect 1542 2913 1548 3978
rect 1660 3016 1666 4085
rect 1700 3016 1706 4085
rect 1792 4096 1892 4098
rect 1792 4044 1816 4096
rect 1868 4044 1892 4096
rect 1792 4032 1892 4044
rect 1792 3980 1816 4032
rect 1868 3980 1892 4032
rect 1792 3978 1892 3980
rect 1976 4085 2022 4097
rect 1516 2909 1548 2913
rect 1502 2897 1548 2909
rect 1632 3014 1732 3016
rect 1632 2962 1656 3014
rect 1708 2962 1732 3014
rect 1632 2950 1732 2962
rect 1632 2898 1656 2950
rect 1708 2898 1732 2950
rect 1632 2896 1732 2898
rect 1818 2909 1824 3978
rect 1858 2909 1864 3978
rect 1976 3016 1982 4085
rect 2016 3016 2022 4085
rect 2108 4096 2208 4098
rect 2108 4044 2132 4096
rect 2184 4044 2208 4096
rect 2108 4032 2208 4044
rect 2108 3980 2132 4032
rect 2184 3980 2208 4032
rect 2108 3978 2208 3980
rect 2292 4085 2338 4101
rect 2394 4100 2446 4122
rect 1818 2897 1864 2909
rect 1948 3014 2048 3016
rect 1948 2962 1972 3014
rect 2024 2962 2048 3014
rect 1948 2950 2048 2962
rect 1948 2898 1972 2950
rect 2024 2898 2048 2950
rect 1948 2896 2048 2898
rect 2134 2909 2140 3978
rect 2174 2909 2180 3978
rect 2292 3016 2298 4085
rect 2332 3016 2338 4085
rect 2370 4098 2450 4100
rect 2370 4046 2384 4098
rect 2436 4093 2450 4098
rect 2437 4059 2450 4093
rect 2436 4046 2450 4059
rect 2370 4034 2450 4046
rect 2370 3982 2384 4034
rect 2436 4021 2450 4034
rect 2437 3987 2450 4021
rect 2436 3982 2450 3987
rect 2370 3980 2450 3982
rect 2394 3958 2446 3980
rect 2134 2897 2180 2909
rect 2264 3014 2364 3016
rect 2264 2962 2288 3014
rect 2340 2962 2364 3014
rect 2264 2950 2364 2962
rect 2264 2898 2288 2950
rect 2340 2898 2364 2950
rect 2264 2896 2364 2898
rect -140 2816 142 2850
rect -140 1484 -70 2816
rect 147 2809 2293 2855
rect 80 2719 126 2731
rect 80 1650 86 2719
rect 120 1650 126 2719
rect 212 2730 312 2732
rect 212 2678 236 2730
rect 288 2678 312 2730
rect 212 2666 312 2678
rect 212 2614 236 2666
rect 288 2614 312 2666
rect 212 2612 312 2614
rect 396 2719 442 2735
rect 52 1648 152 1650
rect 52 1596 76 1648
rect 128 1596 152 1648
rect 52 1584 152 1596
rect 52 1532 76 1584
rect 128 1532 152 1584
rect 52 1530 152 1532
rect 238 1543 244 2612
rect 278 1543 284 2612
rect 396 1650 402 2719
rect 436 1650 442 2719
rect 528 2730 628 2732
rect 528 2678 552 2730
rect 604 2678 628 2730
rect 528 2666 628 2678
rect 528 2614 552 2666
rect 604 2614 628 2666
rect 528 2612 628 2614
rect 712 2719 758 2731
rect 238 1531 284 1543
rect 368 1648 468 1650
rect 368 1596 392 1648
rect 444 1596 468 1648
rect 368 1584 468 1596
rect 368 1532 392 1584
rect 444 1532 468 1584
rect 368 1530 468 1532
rect 554 1543 560 2612
rect 594 1547 600 2612
rect 712 1650 718 2719
rect 752 1650 758 2719
rect 844 2730 944 2732
rect 844 2678 868 2730
rect 920 2678 944 2730
rect 844 2666 944 2678
rect 844 2614 868 2666
rect 920 2614 944 2666
rect 844 2612 944 2614
rect 1028 2719 1074 2731
rect 568 1543 600 1547
rect 554 1531 600 1543
rect 684 1648 784 1650
rect 684 1596 708 1648
rect 760 1596 784 1648
rect 684 1584 784 1596
rect 684 1532 708 1584
rect 760 1532 784 1584
rect 684 1530 784 1532
rect 870 1543 876 2612
rect 910 1543 916 2612
rect 1028 1650 1034 2719
rect 1068 1650 1074 2719
rect 1160 2730 1260 2732
rect 1160 2678 1184 2730
rect 1236 2678 1260 2730
rect 1160 2666 1260 2678
rect 1160 2614 1184 2666
rect 1236 2614 1260 2666
rect 1160 2612 1260 2614
rect 1344 2719 1390 2735
rect 870 1531 916 1543
rect 1000 1648 1100 1650
rect 1000 1596 1024 1648
rect 1076 1596 1100 1648
rect 1000 1584 1100 1596
rect 1000 1532 1024 1584
rect 1076 1532 1100 1584
rect 1000 1530 1100 1532
rect 1186 1543 1192 2612
rect 1226 1543 1232 2612
rect 1344 1650 1350 2719
rect 1384 1650 1390 2719
rect 1476 2730 1576 2732
rect 1476 2678 1500 2730
rect 1552 2678 1576 2730
rect 1476 2666 1576 2678
rect 1476 2614 1500 2666
rect 1552 2614 1576 2666
rect 1476 2612 1576 2614
rect 1660 2719 1706 2731
rect 1186 1531 1232 1543
rect 1316 1648 1416 1650
rect 1316 1596 1340 1648
rect 1392 1596 1416 1648
rect 1316 1584 1416 1596
rect 1316 1532 1340 1584
rect 1392 1532 1416 1584
rect 1316 1530 1416 1532
rect 1502 1543 1508 2612
rect 1542 1547 1548 2612
rect 1660 1650 1666 2719
rect 1700 1650 1706 2719
rect 1792 2730 1892 2732
rect 1792 2678 1816 2730
rect 1868 2678 1892 2730
rect 1792 2666 1892 2678
rect 1792 2614 1816 2666
rect 1868 2614 1892 2666
rect 1792 2612 1892 2614
rect 1976 2719 2022 2731
rect 1516 1543 1548 1547
rect 1502 1531 1548 1543
rect 1632 1648 1732 1650
rect 1632 1596 1656 1648
rect 1708 1596 1732 1648
rect 1632 1584 1732 1596
rect 1632 1532 1656 1584
rect 1708 1532 1732 1584
rect 1632 1530 1732 1532
rect 1818 1543 1824 2612
rect 1858 1543 1864 2612
rect 1976 1650 1982 2719
rect 2016 1650 2022 2719
rect 2108 2730 2208 2732
rect 2108 2678 2132 2730
rect 2184 2678 2208 2730
rect 2108 2666 2208 2678
rect 2108 2614 2132 2666
rect 2184 2614 2208 2666
rect 2108 2612 2208 2614
rect 2292 2719 2338 2735
rect 2394 2730 2446 2752
rect 1818 1531 1864 1543
rect 1948 1648 2048 1650
rect 1948 1596 1972 1648
rect 2024 1596 2048 1648
rect 1948 1584 2048 1596
rect 1948 1532 1972 1584
rect 2024 1532 2048 1584
rect 1948 1530 2048 1532
rect 2134 1543 2140 2612
rect 2174 1543 2180 2612
rect 2292 1650 2298 2719
rect 2332 1650 2338 2719
rect 2370 2728 2450 2730
rect 2370 2676 2384 2728
rect 2436 2723 2450 2728
rect 2437 2689 2450 2723
rect 2436 2676 2450 2689
rect 2370 2664 2450 2676
rect 2370 2612 2384 2664
rect 2436 2651 2450 2664
rect 2437 2617 2450 2651
rect 2436 2612 2450 2617
rect 2370 2610 2450 2612
rect 2394 2588 2446 2610
rect 2134 1531 2180 1543
rect 2264 1648 2364 1650
rect 2264 1596 2288 1648
rect 2340 1596 2364 1648
rect 2264 1584 2364 1596
rect 2264 1532 2288 1584
rect 2340 1532 2364 1584
rect 2264 1530 2364 1532
rect -140 1450 142 1484
rect -140 118 -70 1450
rect 147 1444 2293 1490
rect 80 1353 126 1365
rect 80 284 86 1353
rect 120 284 126 1353
rect 212 1364 312 1366
rect 212 1312 236 1364
rect 288 1312 312 1364
rect 212 1300 312 1312
rect 212 1248 236 1300
rect 288 1248 312 1300
rect 212 1246 312 1248
rect 396 1353 442 1369
rect 52 282 152 284
rect 52 230 76 282
rect 128 230 152 282
rect 52 218 152 230
rect 52 166 76 218
rect 128 166 152 218
rect 52 164 152 166
rect 238 177 244 1246
rect 278 177 284 1246
rect 396 284 402 1353
rect 436 284 442 1353
rect 528 1364 628 1366
rect 528 1312 552 1364
rect 604 1312 628 1364
rect 528 1300 628 1312
rect 528 1248 552 1300
rect 604 1248 628 1300
rect 528 1246 628 1248
rect 712 1353 758 1365
rect 238 165 284 177
rect 368 282 468 284
rect 368 230 392 282
rect 444 230 468 282
rect 368 218 468 230
rect 368 166 392 218
rect 444 166 468 218
rect 368 164 468 166
rect 554 177 560 1246
rect 594 181 600 1246
rect 712 284 718 1353
rect 752 284 758 1353
rect 844 1364 944 1366
rect 844 1312 868 1364
rect 920 1312 944 1364
rect 844 1300 944 1312
rect 844 1248 868 1300
rect 920 1248 944 1300
rect 844 1246 944 1248
rect 1028 1353 1074 1365
rect 568 177 600 181
rect 554 165 600 177
rect 684 282 784 284
rect 684 230 708 282
rect 760 230 784 282
rect 684 218 784 230
rect 684 166 708 218
rect 760 166 784 218
rect 684 164 784 166
rect 870 177 876 1246
rect 910 177 916 1246
rect 1028 284 1034 1353
rect 1068 284 1074 1353
rect 1160 1364 1260 1366
rect 1160 1312 1184 1364
rect 1236 1312 1260 1364
rect 1160 1300 1260 1312
rect 1160 1248 1184 1300
rect 1236 1248 1260 1300
rect 1160 1246 1260 1248
rect 1344 1353 1390 1369
rect 870 165 916 177
rect 1000 282 1100 284
rect 1000 230 1024 282
rect 1076 230 1100 282
rect 1000 218 1100 230
rect 1000 166 1024 218
rect 1076 166 1100 218
rect 1000 164 1100 166
rect 1186 177 1192 1246
rect 1226 177 1232 1246
rect 1344 284 1350 1353
rect 1384 284 1390 1353
rect 1476 1364 1576 1366
rect 1476 1312 1500 1364
rect 1552 1312 1576 1364
rect 1476 1300 1576 1312
rect 1476 1248 1500 1300
rect 1552 1248 1576 1300
rect 1476 1246 1576 1248
rect 1660 1353 1706 1365
rect 1186 165 1232 177
rect 1316 282 1416 284
rect 1316 230 1340 282
rect 1392 230 1416 282
rect 1316 218 1416 230
rect 1316 166 1340 218
rect 1392 166 1416 218
rect 1316 164 1416 166
rect 1502 177 1508 1246
rect 1542 181 1548 1246
rect 1660 284 1666 1353
rect 1700 284 1706 1353
rect 1792 1364 1892 1366
rect 1792 1312 1816 1364
rect 1868 1312 1892 1364
rect 1792 1300 1892 1312
rect 1792 1248 1816 1300
rect 1868 1248 1892 1300
rect 1792 1246 1892 1248
rect 1976 1353 2022 1365
rect 1516 177 1548 181
rect 1502 165 1548 177
rect 1632 282 1732 284
rect 1632 230 1656 282
rect 1708 230 1732 282
rect 1632 218 1732 230
rect 1632 166 1656 218
rect 1708 166 1732 218
rect 1632 164 1732 166
rect 1818 177 1824 1246
rect 1858 177 1864 1246
rect 1976 284 1982 1353
rect 2016 284 2022 1353
rect 2108 1364 2208 1366
rect 2108 1312 2132 1364
rect 2184 1312 2208 1364
rect 2108 1300 2208 1312
rect 2108 1248 2132 1300
rect 2184 1248 2208 1300
rect 2108 1246 2208 1248
rect 2292 1353 2338 1369
rect 2394 1363 2446 1392
rect 2394 1360 2403 1363
rect 1818 165 1864 177
rect 1948 282 2048 284
rect 1948 230 1972 282
rect 2024 230 2048 282
rect 1948 218 2048 230
rect 1948 166 1972 218
rect 2024 166 2048 218
rect 1948 164 2048 166
rect 2134 177 2140 1246
rect 2174 177 2180 1246
rect 2292 284 2298 1353
rect 2332 284 2338 1353
rect 2370 1331 2403 1360
rect 2437 1360 2446 1363
rect 2370 1279 2384 1331
rect 2437 1329 2450 1360
rect 2436 1291 2450 1329
rect 2370 1257 2403 1279
rect 2437 1257 2450 1291
rect 2370 1250 2450 1257
rect 2394 1228 2446 1250
rect 2134 165 2180 177
rect 2264 282 2364 284
rect 2264 230 2288 282
rect 2340 230 2364 282
rect 2264 218 2364 230
rect 2264 166 2288 218
rect 2340 166 2364 218
rect 2264 164 2364 166
rect -140 84 142 118
rect -140 80 -70 84
rect 147 79 2293 125
<< via1 >>
rect 236 5408 288 5460
rect 236 5344 288 5396
rect 552 5408 604 5460
rect 552 5344 604 5396
rect 76 4326 128 4378
rect 76 4262 128 4314
rect 392 4326 444 4378
rect 392 4262 444 4314
rect 868 5408 920 5460
rect 868 5344 920 5396
rect 708 4326 760 4378
rect 708 4262 760 4314
rect 1184 5408 1236 5460
rect 1184 5344 1236 5396
rect 1024 4326 1076 4378
rect 1024 4262 1076 4314
rect 1500 5408 1552 5460
rect 1500 5344 1552 5396
rect 1340 4326 1392 4378
rect 1340 4262 1392 4314
rect 1816 5408 1868 5460
rect 1816 5344 1868 5396
rect 1656 4326 1708 4378
rect 1656 4262 1708 4314
rect 2132 5408 2184 5460
rect 2132 5344 2184 5396
rect 1972 4326 2024 4378
rect 1972 4262 2024 4314
rect 2384 5453 2436 5458
rect 2384 5419 2403 5453
rect 2403 5419 2436 5453
rect 2384 5406 2436 5419
rect 2384 5381 2436 5394
rect 2384 5347 2403 5381
rect 2403 5347 2436 5381
rect 2384 5342 2436 5347
rect 2288 4326 2340 4378
rect 2288 4262 2340 4314
rect 236 4044 288 4096
rect 236 3980 288 4032
rect 76 2962 128 3014
rect 76 2898 128 2950
rect 552 4044 604 4096
rect 552 3980 604 4032
rect 392 2962 444 3014
rect 392 2898 444 2950
rect 868 4044 920 4096
rect 868 3980 920 4032
rect 708 2962 760 3014
rect 708 2898 760 2950
rect 1184 4044 1236 4096
rect 1184 3980 1236 4032
rect 1024 2962 1076 3014
rect 1024 2898 1076 2950
rect 1500 4044 1552 4096
rect 1500 3980 1552 4032
rect 1340 2962 1392 3014
rect 1340 2898 1392 2950
rect 1816 4044 1868 4096
rect 1816 3980 1868 4032
rect 1656 2962 1708 3014
rect 1656 2898 1708 2950
rect 2132 4044 2184 4096
rect 2132 3980 2184 4032
rect 1972 2962 2024 3014
rect 1972 2898 2024 2950
rect 2384 4093 2436 4098
rect 2384 4059 2403 4093
rect 2403 4059 2436 4093
rect 2384 4046 2436 4059
rect 2384 4021 2436 4034
rect 2384 3987 2403 4021
rect 2403 3987 2436 4021
rect 2384 3982 2436 3987
rect 2288 2962 2340 3014
rect 2288 2898 2340 2950
rect 236 2678 288 2730
rect 236 2614 288 2666
rect 76 1596 128 1648
rect 76 1532 128 1584
rect 552 2678 604 2730
rect 552 2614 604 2666
rect 392 1596 444 1648
rect 392 1532 444 1584
rect 868 2678 920 2730
rect 868 2614 920 2666
rect 708 1596 760 1648
rect 708 1532 760 1584
rect 1184 2678 1236 2730
rect 1184 2614 1236 2666
rect 1024 1596 1076 1648
rect 1024 1532 1076 1584
rect 1500 2678 1552 2730
rect 1500 2614 1552 2666
rect 1340 1596 1392 1648
rect 1340 1532 1392 1584
rect 1816 2678 1868 2730
rect 1816 2614 1868 2666
rect 1656 1596 1708 1648
rect 1656 1532 1708 1584
rect 2132 2678 2184 2730
rect 2132 2614 2184 2666
rect 1972 1596 2024 1648
rect 1972 1532 2024 1584
rect 2384 2723 2436 2728
rect 2384 2689 2403 2723
rect 2403 2689 2436 2723
rect 2384 2676 2436 2689
rect 2384 2651 2436 2664
rect 2384 2617 2403 2651
rect 2403 2617 2436 2651
rect 2384 2612 2436 2617
rect 2288 1596 2340 1648
rect 2288 1532 2340 1584
rect 236 1312 288 1364
rect 236 1248 288 1300
rect 76 230 128 282
rect 76 166 128 218
rect 552 1312 604 1364
rect 552 1248 604 1300
rect 392 230 444 282
rect 392 166 444 218
rect 868 1312 920 1364
rect 868 1248 920 1300
rect 708 230 760 282
rect 708 166 760 218
rect 1184 1312 1236 1364
rect 1184 1248 1236 1300
rect 1024 230 1076 282
rect 1024 166 1076 218
rect 1500 1312 1552 1364
rect 1500 1248 1552 1300
rect 1340 230 1392 282
rect 1340 166 1392 218
rect 1816 1312 1868 1364
rect 1816 1248 1868 1300
rect 1656 230 1708 282
rect 1656 166 1708 218
rect 2132 1312 2184 1364
rect 2132 1248 2184 1300
rect 1972 230 2024 282
rect 1972 166 2024 218
rect 2384 1329 2403 1331
rect 2403 1329 2436 1331
rect 2384 1291 2436 1329
rect 2384 1279 2403 1291
rect 2403 1279 2436 1291
rect 2288 230 2340 282
rect 2288 166 2340 218
<< metal2 >>
rect 222 5460 2446 5472
rect 222 5408 236 5460
rect 288 5408 552 5460
rect 604 5408 868 5460
rect 920 5438 1184 5460
rect 1236 5438 1500 5460
rect 920 5408 1142 5438
rect 1278 5408 1500 5438
rect 1552 5408 1816 5460
rect 1868 5408 2132 5460
rect 2184 5458 2446 5460
rect 2184 5408 2384 5458
rect 222 5396 1142 5408
rect 1198 5396 1222 5408
rect 1278 5406 2384 5408
rect 2436 5406 2446 5458
rect 1278 5396 2446 5406
rect 222 5344 236 5396
rect 288 5344 552 5396
rect 604 5344 868 5396
rect 920 5382 1142 5396
rect 1278 5382 1500 5396
rect 920 5344 1184 5382
rect 1236 5344 1500 5382
rect 1552 5344 1816 5396
rect 1868 5344 2132 5396
rect 2184 5394 2446 5396
rect 2184 5344 2384 5394
rect 222 5342 2384 5344
rect 2436 5342 2446 5394
rect 222 5332 2446 5342
rect 2380 5330 2440 5332
rect -40 4378 2354 4390
rect -40 4326 76 4378
rect 128 4326 392 4378
rect 444 4326 708 4378
rect 760 4326 1024 4378
rect 1076 4326 1340 4378
rect 1392 4326 1656 4378
rect 1708 4326 1972 4378
rect 2024 4326 2288 4378
rect 2340 4326 2354 4378
rect -40 4314 2354 4326
rect -40 4262 76 4314
rect 128 4262 392 4314
rect 444 4262 708 4314
rect 760 4262 1024 4314
rect 1076 4262 1340 4314
rect 1392 4262 1656 4314
rect 1708 4262 1972 4314
rect 2024 4262 2288 4314
rect 2340 4262 2354 4314
rect -40 4250 2354 4262
rect -40 3026 140 4250
rect 2380 4108 2440 4110
rect 222 4098 2446 4108
rect 222 4096 2384 4098
rect 222 4044 236 4096
rect 288 4044 552 4096
rect 604 4044 868 4096
rect 920 4058 1184 4096
rect 1236 4058 1500 4096
rect 920 4044 1142 4058
rect 1278 4044 1500 4058
rect 1552 4044 1816 4096
rect 1868 4044 2132 4096
rect 2184 4046 2384 4096
rect 2436 4046 2446 4098
rect 2184 4044 2446 4046
rect 222 4032 1142 4044
rect 1198 4032 1222 4044
rect 1278 4034 2446 4044
rect 1278 4032 2384 4034
rect 222 3980 236 4032
rect 288 3980 552 4032
rect 604 3980 868 4032
rect 920 4002 1142 4032
rect 1278 4002 1500 4032
rect 920 3980 1184 4002
rect 1236 3980 1500 4002
rect 1552 3980 1816 4032
rect 1868 3980 2132 4032
rect 2184 3982 2384 4032
rect 2436 3982 2446 4034
rect 2184 3980 2446 3982
rect 222 3970 2446 3980
rect 222 3968 2198 3970
rect -40 3014 2354 3026
rect -40 2962 76 3014
rect 128 2962 392 3014
rect 444 2962 708 3014
rect 760 2962 1024 3014
rect 1076 2962 1340 3014
rect 1392 2962 1656 3014
rect 1708 2962 1972 3014
rect 2024 2962 2288 3014
rect 2340 2962 2354 3014
rect -40 2950 2354 2962
rect -40 2898 76 2950
rect 128 2898 392 2950
rect 444 2898 708 2950
rect 760 2898 1024 2950
rect 1076 2898 1340 2950
rect 1392 2898 1656 2950
rect 1708 2898 1972 2950
rect 2024 2898 2288 2950
rect 2340 2898 2354 2950
rect -40 2886 2354 2898
rect -40 1660 140 2886
rect 222 2740 2198 2742
rect 222 2730 2446 2740
rect 222 2678 236 2730
rect 288 2678 552 2730
rect 604 2678 868 2730
rect 920 2698 1184 2730
rect 1236 2698 1500 2730
rect 920 2678 1142 2698
rect 1278 2678 1500 2698
rect 1552 2678 1816 2730
rect 1868 2678 2132 2730
rect 2184 2728 2446 2730
rect 2184 2678 2384 2728
rect 222 2666 1142 2678
rect 1198 2666 1222 2678
rect 1278 2676 2384 2678
rect 2436 2676 2446 2728
rect 1278 2666 2446 2676
rect 222 2614 236 2666
rect 288 2614 552 2666
rect 604 2614 868 2666
rect 920 2642 1142 2666
rect 1278 2642 1500 2666
rect 920 2614 1184 2642
rect 1236 2614 1500 2642
rect 1552 2614 1816 2666
rect 1868 2614 2132 2666
rect 2184 2664 2446 2666
rect 2184 2614 2384 2664
rect 222 2612 2384 2614
rect 2436 2612 2446 2664
rect 222 2602 2446 2612
rect 2380 2600 2440 2602
rect -40 1648 2354 1660
rect -40 1596 76 1648
rect 128 1596 392 1648
rect 444 1596 708 1648
rect 760 1596 1024 1648
rect 1076 1596 1340 1648
rect 1392 1596 1656 1648
rect 1708 1596 1972 1648
rect 2024 1596 2288 1648
rect 2340 1596 2354 1648
rect -40 1584 2354 1596
rect -40 1532 76 1584
rect 128 1532 392 1584
rect 444 1532 708 1584
rect 760 1532 1024 1584
rect 1076 1532 1340 1584
rect 1392 1532 1656 1584
rect 1708 1532 1972 1584
rect 2024 1532 2288 1584
rect 2340 1532 2354 1584
rect -40 1520 2354 1532
rect -40 294 140 1520
rect 222 1364 2446 1376
rect 222 1312 236 1364
rect 288 1312 552 1364
rect 604 1312 868 1364
rect 920 1328 1184 1364
rect 1236 1328 1500 1364
rect 920 1312 1142 1328
rect 1278 1312 1500 1328
rect 1552 1312 1816 1364
rect 1868 1312 2132 1364
rect 2184 1331 2446 1364
rect 2184 1312 2384 1331
rect 222 1300 1142 1312
rect 1198 1300 1222 1312
rect 1278 1300 2384 1312
rect 222 1248 236 1300
rect 288 1248 552 1300
rect 604 1248 868 1300
rect 920 1272 1142 1300
rect 1278 1272 1500 1300
rect 920 1248 1184 1272
rect 1236 1248 1500 1272
rect 1552 1248 1816 1300
rect 1868 1248 2132 1300
rect 2184 1279 2384 1300
rect 2436 1279 2446 1331
rect 2184 1248 2446 1279
rect 222 1236 2446 1248
rect 1140 1230 1280 1236
rect -40 282 2354 294
rect -40 230 76 282
rect 128 230 392 282
rect 444 230 708 282
rect 760 230 1024 282
rect 1076 230 1340 282
rect 1392 230 1656 282
rect 1708 230 1972 282
rect 2024 230 2288 282
rect 2340 230 2354 282
rect -40 218 2354 230
rect -40 166 76 218
rect 128 166 392 218
rect 444 166 708 218
rect 760 166 1024 218
rect 1076 166 1340 218
rect 1392 166 1656 218
rect 1708 166 1972 218
rect 2024 166 2288 218
rect 2340 166 2354 218
rect -40 154 2354 166
rect -40 150 140 154
<< via2 >>
rect 1142 5408 1184 5438
rect 1184 5408 1198 5438
rect 1222 5408 1236 5438
rect 1236 5408 1278 5438
rect 1142 5396 1198 5408
rect 1222 5396 1278 5408
rect 1142 5382 1184 5396
rect 1184 5382 1198 5396
rect 1222 5382 1236 5396
rect 1236 5382 1278 5396
rect 1142 4044 1184 4058
rect 1184 4044 1198 4058
rect 1222 4044 1236 4058
rect 1236 4044 1278 4058
rect 1142 4032 1198 4044
rect 1222 4032 1278 4044
rect 1142 4002 1184 4032
rect 1184 4002 1198 4032
rect 1222 4002 1236 4032
rect 1236 4002 1278 4032
rect 1142 2678 1184 2698
rect 1184 2678 1198 2698
rect 1222 2678 1236 2698
rect 1236 2678 1278 2698
rect 1142 2666 1198 2678
rect 1222 2666 1278 2678
rect 1142 2642 1184 2666
rect 1184 2642 1198 2666
rect 1222 2642 1236 2666
rect 1236 2642 1278 2666
rect 1142 1312 1184 1328
rect 1184 1312 1198 1328
rect 1222 1312 1236 1328
rect 1236 1312 1278 1328
rect 1142 1300 1198 1312
rect 1222 1300 1278 1312
rect 1142 1272 1184 1300
rect 1184 1272 1198 1300
rect 1222 1272 1236 1300
rect 1236 1272 1278 1300
<< metal3 >>
rect 1130 5438 1290 5650
rect 1130 5382 1142 5438
rect 1198 5382 1222 5438
rect 1278 5382 1290 5438
rect 1130 4058 1290 5382
rect 1130 4002 1142 4058
rect 1198 4002 1222 4058
rect 1278 4002 1290 4058
rect 1130 2698 1290 4002
rect 1130 2642 1142 2698
rect 1198 2642 1222 2698
rect 1278 2642 1290 2698
rect 1130 1328 1290 2642
rect 1130 1272 1142 1328
rect 1198 1272 1222 1328
rect 1278 1272 1290 1328
rect 1130 1235 1290 1272
use sky130_fd_pr__pfet_01v8_lvt_D74VRS  sky130_fd_pr__pfet_01v8_lvt_D74VRS_0
timestamp 1663011646
transform 1 0 1209 0 1 2778
box -1273 -2831 1273 2831
<< end >>
