magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -159 -111 -97 -105
rect -31 -111 31 -105
rect 97 -111 159 -105
rect -159 -145 -145 -111
rect -31 -145 -17 -111
rect 97 -145 111 -111
rect -159 -151 -97 -145
rect -31 -151 31 -145
rect 97 -151 159 -145
<< nwell >>
rect -359 -284 359 284
<< pmoslvt >>
rect -163 -64 -93 136
rect -35 -64 35 136
rect 93 -64 163 136
<< pdiff >>
rect -221 121 -163 136
rect -221 87 -209 121
rect -175 87 -163 121
rect -221 53 -163 87
rect -221 19 -209 53
rect -175 19 -163 53
rect -221 -15 -163 19
rect -221 -49 -209 -15
rect -175 -49 -163 -15
rect -221 -64 -163 -49
rect -93 121 -35 136
rect -93 87 -81 121
rect -47 87 -35 121
rect -93 53 -35 87
rect -93 19 -81 53
rect -47 19 -35 53
rect -93 -15 -35 19
rect -93 -49 -81 -15
rect -47 -49 -35 -15
rect -93 -64 -35 -49
rect 35 121 93 136
rect 35 87 47 121
rect 81 87 93 121
rect 35 53 93 87
rect 35 19 47 53
rect 81 19 93 53
rect 35 -15 93 19
rect 35 -49 47 -15
rect 81 -49 93 -15
rect 35 -64 93 -49
rect 163 121 221 136
rect 163 87 175 121
rect 209 87 221 121
rect 163 53 221 87
rect 163 19 175 53
rect 209 19 221 53
rect 163 -15 221 19
rect 163 -49 175 -15
rect 209 -49 221 -15
rect 163 -64 221 -49
<< pdiffc >>
rect -209 87 -175 121
rect -209 19 -175 53
rect -209 -49 -175 -15
rect -81 87 -47 121
rect -81 19 -47 53
rect -81 -49 -47 -15
rect 47 87 81 121
rect 47 19 81 53
rect 47 -49 81 -15
rect 175 87 209 121
rect 175 19 209 53
rect 175 -49 209 -15
<< nsubdiff >>
rect -323 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 323 248
rect -323 119 -289 214
rect -323 51 -289 85
rect -323 -17 -289 17
rect -323 -85 -289 -51
rect 289 119 323 214
rect 289 51 323 85
rect 289 -17 323 17
rect -323 -214 -289 -119
rect 289 -85 323 -51
rect 289 -214 323 -119
rect -323 -248 -221 -214
rect -187 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 187 -214
rect 221 -248 323 -214
<< nsubdiffcont >>
rect -221 214 -187 248
rect -153 214 -119 248
rect -85 214 -51 248
rect -17 214 17 248
rect 51 214 85 248
rect 119 214 153 248
rect 187 214 221 248
rect -323 85 -289 119
rect -323 17 -289 51
rect -323 -51 -289 -17
rect 289 85 323 119
rect 289 17 323 51
rect 289 -51 323 -17
rect -323 -119 -289 -85
rect 289 -119 323 -85
rect -221 -248 -187 -214
rect -153 -248 -119 -214
rect -85 -248 -51 -214
rect -17 -248 17 -214
rect 51 -248 85 -214
rect 119 -248 153 -214
rect 187 -248 221 -214
<< poly >>
rect -163 136 -93 162
rect -35 136 35 162
rect 93 136 163 162
rect -163 -111 -93 -64
rect -163 -145 -145 -111
rect -111 -145 -93 -111
rect -163 -161 -93 -145
rect -35 -111 35 -64
rect -35 -145 -17 -111
rect 17 -145 35 -111
rect -35 -161 35 -145
rect 93 -111 163 -64
rect 93 -145 111 -111
rect 145 -145 163 -111
rect 93 -161 163 -145
<< polycont >>
rect -145 -145 -111 -111
rect -17 -145 17 -111
rect 111 -145 145 -111
<< locali >>
rect -323 214 -221 248
rect -187 214 -153 248
rect -119 214 -85 248
rect -51 214 -17 248
rect 17 214 51 248
rect 85 214 119 248
rect 153 214 187 248
rect 221 214 323 248
rect -323 119 -289 214
rect -323 51 -289 85
rect -323 -17 -289 17
rect -323 -85 -289 -51
rect -209 121 -175 140
rect -209 53 -175 55
rect -209 17 -175 19
rect -209 -68 -175 -49
rect -81 121 -47 140
rect -81 53 -47 55
rect -81 17 -47 19
rect -81 -68 -47 -49
rect 47 121 81 140
rect 47 53 81 55
rect 47 17 81 19
rect 47 -68 81 -49
rect 175 121 209 140
rect 175 53 209 55
rect 175 17 209 19
rect 175 -68 209 -49
rect 289 119 323 214
rect 289 51 323 85
rect 289 -17 323 17
rect 289 -85 323 -51
rect -323 -214 -289 -119
rect -163 -145 -145 -111
rect -111 -145 -93 -111
rect -35 -145 -17 -111
rect 17 -145 35 -111
rect 93 -145 111 -111
rect 145 -145 163 -111
rect 289 -214 323 -119
rect -323 -248 -221 -214
rect -187 -248 -153 -214
rect -119 -248 -85 -214
rect -51 -248 -17 -214
rect 17 -248 51 -214
rect 85 -248 119 -214
rect 153 -248 187 -214
rect 221 -248 323 -214
<< viali >>
rect -209 87 -175 89
rect -209 55 -175 87
rect -209 -15 -175 17
rect -209 -17 -175 -15
rect -81 87 -47 89
rect -81 55 -47 87
rect -81 -15 -47 17
rect -81 -17 -47 -15
rect 47 87 81 89
rect 47 55 81 87
rect 47 -15 81 17
rect 47 -17 81 -15
rect 175 87 209 89
rect 175 55 209 87
rect 175 -15 209 17
rect 175 -17 209 -15
rect -145 -145 -111 -111
rect -17 -145 17 -111
rect 111 -145 145 -111
<< metal1 >>
rect -215 89 -169 136
rect -215 55 -209 89
rect -175 55 -169 89
rect -215 17 -169 55
rect -215 -17 -209 17
rect -175 -17 -169 17
rect -215 -64 -169 -17
rect -87 89 -41 136
rect -87 55 -81 89
rect -47 55 -41 89
rect -87 17 -41 55
rect -87 -17 -81 17
rect -47 -17 -41 17
rect -87 -64 -41 -17
rect 41 89 87 136
rect 41 55 47 89
rect 81 55 87 89
rect 41 17 87 55
rect 41 -17 47 17
rect 81 -17 87 17
rect 41 -64 87 -17
rect 169 89 215 136
rect 169 55 175 89
rect 209 55 215 89
rect 169 17 215 55
rect 169 -17 175 17
rect 209 -17 215 17
rect 169 -64 215 -17
rect -159 -111 -97 -105
rect -159 -145 -145 -111
rect -111 -145 -97 -111
rect -159 -151 -97 -145
rect -31 -111 31 -105
rect -31 -145 -17 -111
rect 17 -145 31 -111
rect -31 -151 31 -145
rect 97 -111 159 -105
rect 97 -145 111 -111
rect 145 -145 159 -111
rect 97 -151 159 -145
<< properties >>
string FIXED_BBOX -306 -231 306 231
<< end >>
