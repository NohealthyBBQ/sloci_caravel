magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -571 -507 571 445
<< nmoslvt >>
rect -487 -481 -287 419
rect -229 -481 -29 419
rect 29 -481 229 419
rect 287 -481 487 419
<< ndiff >>
rect -545 394 -487 419
rect -545 360 -533 394
rect -499 360 -487 394
rect -545 326 -487 360
rect -545 292 -533 326
rect -499 292 -487 326
rect -545 258 -487 292
rect -545 224 -533 258
rect -499 224 -487 258
rect -545 190 -487 224
rect -545 156 -533 190
rect -499 156 -487 190
rect -545 122 -487 156
rect -545 88 -533 122
rect -499 88 -487 122
rect -545 54 -487 88
rect -545 20 -533 54
rect -499 20 -487 54
rect -545 -14 -487 20
rect -545 -48 -533 -14
rect -499 -48 -487 -14
rect -545 -82 -487 -48
rect -545 -116 -533 -82
rect -499 -116 -487 -82
rect -545 -150 -487 -116
rect -545 -184 -533 -150
rect -499 -184 -487 -150
rect -545 -218 -487 -184
rect -545 -252 -533 -218
rect -499 -252 -487 -218
rect -545 -286 -487 -252
rect -545 -320 -533 -286
rect -499 -320 -487 -286
rect -545 -354 -487 -320
rect -545 -388 -533 -354
rect -499 -388 -487 -354
rect -545 -422 -487 -388
rect -545 -456 -533 -422
rect -499 -456 -487 -422
rect -545 -481 -487 -456
rect -287 394 -229 419
rect -287 360 -275 394
rect -241 360 -229 394
rect -287 326 -229 360
rect -287 292 -275 326
rect -241 292 -229 326
rect -287 258 -229 292
rect -287 224 -275 258
rect -241 224 -229 258
rect -287 190 -229 224
rect -287 156 -275 190
rect -241 156 -229 190
rect -287 122 -229 156
rect -287 88 -275 122
rect -241 88 -229 122
rect -287 54 -229 88
rect -287 20 -275 54
rect -241 20 -229 54
rect -287 -14 -229 20
rect -287 -48 -275 -14
rect -241 -48 -229 -14
rect -287 -82 -229 -48
rect -287 -116 -275 -82
rect -241 -116 -229 -82
rect -287 -150 -229 -116
rect -287 -184 -275 -150
rect -241 -184 -229 -150
rect -287 -218 -229 -184
rect -287 -252 -275 -218
rect -241 -252 -229 -218
rect -287 -286 -229 -252
rect -287 -320 -275 -286
rect -241 -320 -229 -286
rect -287 -354 -229 -320
rect -287 -388 -275 -354
rect -241 -388 -229 -354
rect -287 -422 -229 -388
rect -287 -456 -275 -422
rect -241 -456 -229 -422
rect -287 -481 -229 -456
rect -29 394 29 419
rect -29 360 -17 394
rect 17 360 29 394
rect -29 326 29 360
rect -29 292 -17 326
rect 17 292 29 326
rect -29 258 29 292
rect -29 224 -17 258
rect 17 224 29 258
rect -29 190 29 224
rect -29 156 -17 190
rect 17 156 29 190
rect -29 122 29 156
rect -29 88 -17 122
rect 17 88 29 122
rect -29 54 29 88
rect -29 20 -17 54
rect 17 20 29 54
rect -29 -14 29 20
rect -29 -48 -17 -14
rect 17 -48 29 -14
rect -29 -82 29 -48
rect -29 -116 -17 -82
rect 17 -116 29 -82
rect -29 -150 29 -116
rect -29 -184 -17 -150
rect 17 -184 29 -150
rect -29 -218 29 -184
rect -29 -252 -17 -218
rect 17 -252 29 -218
rect -29 -286 29 -252
rect -29 -320 -17 -286
rect 17 -320 29 -286
rect -29 -354 29 -320
rect -29 -388 -17 -354
rect 17 -388 29 -354
rect -29 -422 29 -388
rect -29 -456 -17 -422
rect 17 -456 29 -422
rect -29 -481 29 -456
rect 229 394 287 419
rect 229 360 241 394
rect 275 360 287 394
rect 229 326 287 360
rect 229 292 241 326
rect 275 292 287 326
rect 229 258 287 292
rect 229 224 241 258
rect 275 224 287 258
rect 229 190 287 224
rect 229 156 241 190
rect 275 156 287 190
rect 229 122 287 156
rect 229 88 241 122
rect 275 88 287 122
rect 229 54 287 88
rect 229 20 241 54
rect 275 20 287 54
rect 229 -14 287 20
rect 229 -48 241 -14
rect 275 -48 287 -14
rect 229 -82 287 -48
rect 229 -116 241 -82
rect 275 -116 287 -82
rect 229 -150 287 -116
rect 229 -184 241 -150
rect 275 -184 287 -150
rect 229 -218 287 -184
rect 229 -252 241 -218
rect 275 -252 287 -218
rect 229 -286 287 -252
rect 229 -320 241 -286
rect 275 -320 287 -286
rect 229 -354 287 -320
rect 229 -388 241 -354
rect 275 -388 287 -354
rect 229 -422 287 -388
rect 229 -456 241 -422
rect 275 -456 287 -422
rect 229 -481 287 -456
rect 487 394 545 419
rect 487 360 499 394
rect 533 360 545 394
rect 487 326 545 360
rect 487 292 499 326
rect 533 292 545 326
rect 487 258 545 292
rect 487 224 499 258
rect 533 224 545 258
rect 487 190 545 224
rect 487 156 499 190
rect 533 156 545 190
rect 487 122 545 156
rect 487 88 499 122
rect 533 88 545 122
rect 487 54 545 88
rect 487 20 499 54
rect 533 20 545 54
rect 487 -14 545 20
rect 487 -48 499 -14
rect 533 -48 545 -14
rect 487 -82 545 -48
rect 487 -116 499 -82
rect 533 -116 545 -82
rect 487 -150 545 -116
rect 487 -184 499 -150
rect 533 -184 545 -150
rect 487 -218 545 -184
rect 487 -252 499 -218
rect 533 -252 545 -218
rect 487 -286 545 -252
rect 487 -320 499 -286
rect 533 -320 545 -286
rect 487 -354 545 -320
rect 487 -388 499 -354
rect 533 -388 545 -354
rect 487 -422 545 -388
rect 487 -456 499 -422
rect 533 -456 545 -422
rect 487 -481 545 -456
<< ndiffc >>
rect -533 360 -499 394
rect -533 292 -499 326
rect -533 224 -499 258
rect -533 156 -499 190
rect -533 88 -499 122
rect -533 20 -499 54
rect -533 -48 -499 -14
rect -533 -116 -499 -82
rect -533 -184 -499 -150
rect -533 -252 -499 -218
rect -533 -320 -499 -286
rect -533 -388 -499 -354
rect -533 -456 -499 -422
rect -275 360 -241 394
rect -275 292 -241 326
rect -275 224 -241 258
rect -275 156 -241 190
rect -275 88 -241 122
rect -275 20 -241 54
rect -275 -48 -241 -14
rect -275 -116 -241 -82
rect -275 -184 -241 -150
rect -275 -252 -241 -218
rect -275 -320 -241 -286
rect -275 -388 -241 -354
rect -275 -456 -241 -422
rect -17 360 17 394
rect -17 292 17 326
rect -17 224 17 258
rect -17 156 17 190
rect -17 88 17 122
rect -17 20 17 54
rect -17 -48 17 -14
rect -17 -116 17 -82
rect -17 -184 17 -150
rect -17 -252 17 -218
rect -17 -320 17 -286
rect -17 -388 17 -354
rect -17 -456 17 -422
rect 241 360 275 394
rect 241 292 275 326
rect 241 224 275 258
rect 241 156 275 190
rect 241 88 275 122
rect 241 20 275 54
rect 241 -48 275 -14
rect 241 -116 275 -82
rect 241 -184 275 -150
rect 241 -252 275 -218
rect 241 -320 275 -286
rect 241 -388 275 -354
rect 241 -456 275 -422
rect 499 360 533 394
rect 499 292 533 326
rect 499 224 533 258
rect 499 156 533 190
rect 499 88 533 122
rect 499 20 533 54
rect 499 -48 533 -14
rect 499 -116 533 -82
rect 499 -184 533 -150
rect 499 -252 533 -218
rect 499 -320 533 -286
rect 499 -388 533 -354
rect 499 -456 533 -422
<< poly >>
rect -487 491 -287 507
rect -487 457 -438 491
rect -404 457 -370 491
rect -336 457 -287 491
rect -487 419 -287 457
rect -229 491 -29 507
rect -229 457 -180 491
rect -146 457 -112 491
rect -78 457 -29 491
rect -229 419 -29 457
rect 29 491 229 507
rect 29 457 78 491
rect 112 457 146 491
rect 180 457 229 491
rect 29 419 229 457
rect 287 491 487 507
rect 287 457 336 491
rect 370 457 404 491
rect 438 457 487 491
rect 287 419 487 457
rect -487 -507 -287 -481
rect -229 -507 -29 -481
rect 29 -507 229 -481
rect 287 -507 487 -481
<< polycont >>
rect -438 457 -404 491
rect -370 457 -336 491
rect -180 457 -146 491
rect -112 457 -78 491
rect 78 457 112 491
rect 146 457 180 491
rect 336 457 370 491
rect 404 457 438 491
<< locali >>
rect -487 457 -440 491
rect -404 457 -370 491
rect -334 457 -287 491
rect -229 457 -182 491
rect -146 457 -112 491
rect -76 457 -29 491
rect 29 457 76 491
rect 112 457 146 491
rect 182 457 229 491
rect 287 457 334 491
rect 370 457 404 491
rect 440 457 487 491
rect -533 394 -499 423
rect -533 326 -499 348
rect -533 258 -499 276
rect -533 190 -499 204
rect -533 122 -499 132
rect -533 54 -499 60
rect -533 -14 -499 -12
rect -533 -50 -499 -48
rect -533 -122 -499 -116
rect -533 -194 -499 -184
rect -533 -266 -499 -252
rect -533 -338 -499 -320
rect -533 -410 -499 -388
rect -533 -485 -499 -456
rect -275 394 -241 423
rect -275 326 -241 348
rect -275 258 -241 276
rect -275 190 -241 204
rect -275 122 -241 132
rect -275 54 -241 60
rect -275 -14 -241 -12
rect -275 -50 -241 -48
rect -275 -122 -241 -116
rect -275 -194 -241 -184
rect -275 -266 -241 -252
rect -275 -338 -241 -320
rect -275 -410 -241 -388
rect -275 -485 -241 -456
rect -17 394 17 423
rect -17 326 17 348
rect -17 258 17 276
rect -17 190 17 204
rect -17 122 17 132
rect -17 54 17 60
rect -17 -14 17 -12
rect -17 -50 17 -48
rect -17 -122 17 -116
rect -17 -194 17 -184
rect -17 -266 17 -252
rect -17 -338 17 -320
rect -17 -410 17 -388
rect -17 -485 17 -456
rect 241 394 275 423
rect 241 326 275 348
rect 241 258 275 276
rect 241 190 275 204
rect 241 122 275 132
rect 241 54 275 60
rect 241 -14 275 -12
rect 241 -50 275 -48
rect 241 -122 275 -116
rect 241 -194 275 -184
rect 241 -266 275 -252
rect 241 -338 275 -320
rect 241 -410 275 -388
rect 241 -485 275 -456
rect 499 394 533 423
rect 499 326 533 348
rect 499 258 533 276
rect 499 190 533 204
rect 499 122 533 132
rect 499 54 533 60
rect 499 -14 533 -12
rect 499 -50 533 -48
rect 499 -122 533 -116
rect 499 -194 533 -184
rect 499 -266 533 -252
rect 499 -338 533 -320
rect 499 -410 533 -388
rect 499 -485 533 -456
<< viali >>
rect -440 457 -438 491
rect -438 457 -406 491
rect -368 457 -336 491
rect -336 457 -334 491
rect -182 457 -180 491
rect -180 457 -148 491
rect -110 457 -78 491
rect -78 457 -76 491
rect 76 457 78 491
rect 78 457 110 491
rect 148 457 180 491
rect 180 457 182 491
rect 334 457 336 491
rect 336 457 368 491
rect 406 457 438 491
rect 438 457 440 491
rect -533 360 -499 382
rect -533 348 -499 360
rect -533 292 -499 310
rect -533 276 -499 292
rect -533 224 -499 238
rect -533 204 -499 224
rect -533 156 -499 166
rect -533 132 -499 156
rect -533 88 -499 94
rect -533 60 -499 88
rect -533 20 -499 22
rect -533 -12 -499 20
rect -533 -82 -499 -50
rect -533 -84 -499 -82
rect -533 -150 -499 -122
rect -533 -156 -499 -150
rect -533 -218 -499 -194
rect -533 -228 -499 -218
rect -533 -286 -499 -266
rect -533 -300 -499 -286
rect -533 -354 -499 -338
rect -533 -372 -499 -354
rect -533 -422 -499 -410
rect -533 -444 -499 -422
rect -275 360 -241 382
rect -275 348 -241 360
rect -275 292 -241 310
rect -275 276 -241 292
rect -275 224 -241 238
rect -275 204 -241 224
rect -275 156 -241 166
rect -275 132 -241 156
rect -275 88 -241 94
rect -275 60 -241 88
rect -275 20 -241 22
rect -275 -12 -241 20
rect -275 -82 -241 -50
rect -275 -84 -241 -82
rect -275 -150 -241 -122
rect -275 -156 -241 -150
rect -275 -218 -241 -194
rect -275 -228 -241 -218
rect -275 -286 -241 -266
rect -275 -300 -241 -286
rect -275 -354 -241 -338
rect -275 -372 -241 -354
rect -275 -422 -241 -410
rect -275 -444 -241 -422
rect -17 360 17 382
rect -17 348 17 360
rect -17 292 17 310
rect -17 276 17 292
rect -17 224 17 238
rect -17 204 17 224
rect -17 156 17 166
rect -17 132 17 156
rect -17 88 17 94
rect -17 60 17 88
rect -17 20 17 22
rect -17 -12 17 20
rect -17 -82 17 -50
rect -17 -84 17 -82
rect -17 -150 17 -122
rect -17 -156 17 -150
rect -17 -218 17 -194
rect -17 -228 17 -218
rect -17 -286 17 -266
rect -17 -300 17 -286
rect -17 -354 17 -338
rect -17 -372 17 -354
rect -17 -422 17 -410
rect -17 -444 17 -422
rect 241 360 275 382
rect 241 348 275 360
rect 241 292 275 310
rect 241 276 275 292
rect 241 224 275 238
rect 241 204 275 224
rect 241 156 275 166
rect 241 132 275 156
rect 241 88 275 94
rect 241 60 275 88
rect 241 20 275 22
rect 241 -12 275 20
rect 241 -82 275 -50
rect 241 -84 275 -82
rect 241 -150 275 -122
rect 241 -156 275 -150
rect 241 -218 275 -194
rect 241 -228 275 -218
rect 241 -286 275 -266
rect 241 -300 275 -286
rect 241 -354 275 -338
rect 241 -372 275 -354
rect 241 -422 275 -410
rect 241 -444 275 -422
rect 499 360 533 382
rect 499 348 533 360
rect 499 292 533 310
rect 499 276 533 292
rect 499 224 533 238
rect 499 204 533 224
rect 499 156 533 166
rect 499 132 533 156
rect 499 88 533 94
rect 499 60 533 88
rect 499 20 533 22
rect 499 -12 533 20
rect 499 -82 533 -50
rect 499 -84 533 -82
rect 499 -150 533 -122
rect 499 -156 533 -150
rect 499 -218 533 -194
rect 499 -228 533 -218
rect 499 -286 533 -266
rect 499 -300 533 -286
rect 499 -354 533 -338
rect 499 -372 533 -354
rect 499 -422 533 -410
rect 499 -444 533 -422
<< metal1 >>
rect -483 491 -291 497
rect -483 457 -440 491
rect -406 457 -368 491
rect -334 457 -291 491
rect -483 451 -291 457
rect -225 491 -33 497
rect -225 457 -182 491
rect -148 457 -110 491
rect -76 457 -33 491
rect -225 451 -33 457
rect 33 491 225 497
rect 33 457 76 491
rect 110 457 148 491
rect 182 457 225 491
rect 33 451 225 457
rect 291 491 483 497
rect 291 457 334 491
rect 368 457 406 491
rect 440 457 483 491
rect 291 451 483 457
rect -539 382 -493 419
rect -539 348 -533 382
rect -499 348 -493 382
rect -539 310 -493 348
rect -539 276 -533 310
rect -499 276 -493 310
rect -539 238 -493 276
rect -539 204 -533 238
rect -499 204 -493 238
rect -539 166 -493 204
rect -539 132 -533 166
rect -499 132 -493 166
rect -539 94 -493 132
rect -539 60 -533 94
rect -499 60 -493 94
rect -539 22 -493 60
rect -539 -12 -533 22
rect -499 -12 -493 22
rect -539 -50 -493 -12
rect -539 -84 -533 -50
rect -499 -84 -493 -50
rect -539 -122 -493 -84
rect -539 -156 -533 -122
rect -499 -156 -493 -122
rect -539 -194 -493 -156
rect -539 -228 -533 -194
rect -499 -228 -493 -194
rect -539 -266 -493 -228
rect -539 -300 -533 -266
rect -499 -300 -493 -266
rect -539 -338 -493 -300
rect -539 -372 -533 -338
rect -499 -372 -493 -338
rect -539 -410 -493 -372
rect -539 -444 -533 -410
rect -499 -444 -493 -410
rect -539 -481 -493 -444
rect -281 382 -235 419
rect -281 348 -275 382
rect -241 348 -235 382
rect -281 310 -235 348
rect -281 276 -275 310
rect -241 276 -235 310
rect -281 238 -235 276
rect -281 204 -275 238
rect -241 204 -235 238
rect -281 166 -235 204
rect -281 132 -275 166
rect -241 132 -235 166
rect -281 94 -235 132
rect -281 60 -275 94
rect -241 60 -235 94
rect -281 22 -235 60
rect -281 -12 -275 22
rect -241 -12 -235 22
rect -281 -50 -235 -12
rect -281 -84 -275 -50
rect -241 -84 -235 -50
rect -281 -122 -235 -84
rect -281 -156 -275 -122
rect -241 -156 -235 -122
rect -281 -194 -235 -156
rect -281 -228 -275 -194
rect -241 -228 -235 -194
rect -281 -266 -235 -228
rect -281 -300 -275 -266
rect -241 -300 -235 -266
rect -281 -338 -235 -300
rect -281 -372 -275 -338
rect -241 -372 -235 -338
rect -281 -410 -235 -372
rect -281 -444 -275 -410
rect -241 -444 -235 -410
rect -281 -481 -235 -444
rect -23 382 23 419
rect -23 348 -17 382
rect 17 348 23 382
rect -23 310 23 348
rect -23 276 -17 310
rect 17 276 23 310
rect -23 238 23 276
rect -23 204 -17 238
rect 17 204 23 238
rect -23 166 23 204
rect -23 132 -17 166
rect 17 132 23 166
rect -23 94 23 132
rect -23 60 -17 94
rect 17 60 23 94
rect -23 22 23 60
rect -23 -12 -17 22
rect 17 -12 23 22
rect -23 -50 23 -12
rect -23 -84 -17 -50
rect 17 -84 23 -50
rect -23 -122 23 -84
rect -23 -156 -17 -122
rect 17 -156 23 -122
rect -23 -194 23 -156
rect -23 -228 -17 -194
rect 17 -228 23 -194
rect -23 -266 23 -228
rect -23 -300 -17 -266
rect 17 -300 23 -266
rect -23 -338 23 -300
rect -23 -372 -17 -338
rect 17 -372 23 -338
rect -23 -410 23 -372
rect -23 -444 -17 -410
rect 17 -444 23 -410
rect -23 -481 23 -444
rect 235 382 281 419
rect 235 348 241 382
rect 275 348 281 382
rect 235 310 281 348
rect 235 276 241 310
rect 275 276 281 310
rect 235 238 281 276
rect 235 204 241 238
rect 275 204 281 238
rect 235 166 281 204
rect 235 132 241 166
rect 275 132 281 166
rect 235 94 281 132
rect 235 60 241 94
rect 275 60 281 94
rect 235 22 281 60
rect 235 -12 241 22
rect 275 -12 281 22
rect 235 -50 281 -12
rect 235 -84 241 -50
rect 275 -84 281 -50
rect 235 -122 281 -84
rect 235 -156 241 -122
rect 275 -156 281 -122
rect 235 -194 281 -156
rect 235 -228 241 -194
rect 275 -228 281 -194
rect 235 -266 281 -228
rect 235 -300 241 -266
rect 275 -300 281 -266
rect 235 -338 281 -300
rect 235 -372 241 -338
rect 275 -372 281 -338
rect 235 -410 281 -372
rect 235 -444 241 -410
rect 275 -444 281 -410
rect 235 -481 281 -444
rect 493 382 539 419
rect 493 348 499 382
rect 533 348 539 382
rect 493 310 539 348
rect 493 276 499 310
rect 533 276 539 310
rect 493 238 539 276
rect 493 204 499 238
rect 533 204 539 238
rect 493 166 539 204
rect 493 132 499 166
rect 533 132 539 166
rect 493 94 539 132
rect 493 60 499 94
rect 533 60 539 94
rect 493 22 539 60
rect 493 -12 499 22
rect 533 -12 539 22
rect 493 -50 539 -12
rect 493 -84 499 -50
rect 533 -84 539 -50
rect 493 -122 539 -84
rect 493 -156 499 -122
rect 533 -156 539 -122
rect 493 -194 539 -156
rect 493 -228 499 -194
rect 533 -228 539 -194
rect 493 -266 539 -228
rect 493 -300 499 -266
rect 533 -300 539 -266
rect 493 -338 539 -300
rect 493 -372 499 -338
rect 533 -372 539 -338
rect 493 -410 539 -372
rect 493 -444 499 -410
rect 533 -444 539 -410
rect 493 -481 539 -444
<< end >>
