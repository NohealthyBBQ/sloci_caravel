magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -220 -1060 4440 720
<< nsubdiff >>
rect -140 627 4360 640
rect -140 593 537 627
rect 571 593 605 627
rect 639 593 673 627
rect 707 593 741 627
rect 775 593 809 627
rect 843 593 1317 627
rect 1351 593 1385 627
rect 1419 593 1453 627
rect 1487 593 1521 627
rect 1555 593 1589 627
rect 1623 593 2597 627
rect 2631 593 2665 627
rect 2699 593 2733 627
rect 2767 593 2801 627
rect 2835 593 2869 627
rect 2903 593 3377 627
rect 3411 593 3445 627
rect 3479 593 3513 627
rect 3547 593 3581 627
rect 3615 593 3649 627
rect 3683 593 4360 627
rect -140 580 4360 593
rect -140 447 -80 580
rect -140 413 -127 447
rect -93 413 -80 447
rect -140 379 -80 413
rect -140 345 -127 379
rect -93 345 -80 379
rect -140 311 -80 345
rect -140 277 -127 311
rect -93 277 -80 311
rect -140 243 -80 277
rect -140 209 -127 243
rect -93 209 -80 243
rect -140 175 -80 209
rect -140 141 -127 175
rect -93 141 -80 175
rect -140 107 -80 141
rect -140 73 -127 107
rect -93 73 -80 107
rect -140 -140 -80 73
rect 4300 447 4360 580
rect 4300 413 4313 447
rect 4347 413 4360 447
rect 4300 379 4360 413
rect 4300 345 4313 379
rect 4347 345 4360 379
rect 4300 311 4360 345
rect 4300 277 4313 311
rect 4347 277 4360 311
rect 4300 243 4360 277
rect 4300 209 4313 243
rect 4347 209 4360 243
rect 4300 175 4360 209
rect 4300 141 4313 175
rect 4347 141 4360 175
rect 4300 107 4360 141
rect 4300 73 4313 107
rect 4347 73 4360 107
rect 4300 -140 4360 73
rect -140 -153 4360 -140
rect -140 -187 537 -153
rect 571 -187 605 -153
rect 639 -187 673 -153
rect 707 -187 741 -153
rect 775 -187 809 -153
rect 843 -187 1317 -153
rect 1351 -187 1385 -153
rect 1419 -187 1453 -153
rect 1487 -187 1521 -153
rect 1555 -187 1589 -153
rect 1623 -187 2597 -153
rect 2631 -187 2665 -153
rect 2699 -187 2733 -153
rect 2767 -187 2801 -153
rect 2835 -187 2869 -153
rect 2903 -187 3377 -153
rect 3411 -187 3445 -153
rect 3479 -187 3513 -153
rect 3547 -187 3581 -153
rect 3615 -187 3649 -153
rect 3683 -187 4360 -153
rect -140 -200 4360 -187
rect -140 -413 -80 -200
rect -140 -447 -127 -413
rect -93 -447 -80 -413
rect -140 -481 -80 -447
rect -140 -515 -127 -481
rect -93 -515 -80 -481
rect -140 -549 -80 -515
rect -140 -583 -127 -549
rect -93 -583 -80 -549
rect -140 -617 -80 -583
rect -140 -651 -127 -617
rect -93 -651 -80 -617
rect -140 -685 -80 -651
rect -140 -719 -127 -685
rect -93 -719 -80 -685
rect -140 -753 -80 -719
rect -140 -787 -127 -753
rect -93 -787 -80 -753
rect -140 -920 -80 -787
rect 4300 -413 4360 -200
rect 4300 -447 4313 -413
rect 4347 -447 4360 -413
rect 4300 -481 4360 -447
rect 4300 -515 4313 -481
rect 4347 -515 4360 -481
rect 4300 -549 4360 -515
rect 4300 -583 4313 -549
rect 4347 -583 4360 -549
rect 4300 -617 4360 -583
rect 4300 -651 4313 -617
rect 4347 -651 4360 -617
rect 4300 -685 4360 -651
rect 4300 -719 4313 -685
rect 4347 -719 4360 -685
rect 4300 -753 4360 -719
rect 4300 -787 4313 -753
rect 4347 -787 4360 -753
rect 4300 -920 4360 -787
rect -140 -933 4360 -920
rect -140 -967 537 -933
rect 571 -967 605 -933
rect 639 -967 673 -933
rect 707 -967 741 -933
rect 775 -967 809 -933
rect 843 -967 1317 -933
rect 1351 -967 1385 -933
rect 1419 -967 1453 -933
rect 1487 -967 1521 -933
rect 1555 -967 1589 -933
rect 1623 -967 2597 -933
rect 2631 -967 2665 -933
rect 2699 -967 2733 -933
rect 2767 -967 2801 -933
rect 2835 -967 2869 -933
rect 2903 -967 3377 -933
rect 3411 -967 3445 -933
rect 3479 -967 3513 -933
rect 3547 -967 3581 -933
rect 3615 -967 3649 -933
rect 3683 -967 4360 -933
rect -140 -980 4360 -967
<< nsubdiffcont >>
rect 537 593 571 627
rect 605 593 639 627
rect 673 593 707 627
rect 741 593 775 627
rect 809 593 843 627
rect 1317 593 1351 627
rect 1385 593 1419 627
rect 1453 593 1487 627
rect 1521 593 1555 627
rect 1589 593 1623 627
rect 2597 593 2631 627
rect 2665 593 2699 627
rect 2733 593 2767 627
rect 2801 593 2835 627
rect 2869 593 2903 627
rect 3377 593 3411 627
rect 3445 593 3479 627
rect 3513 593 3547 627
rect 3581 593 3615 627
rect 3649 593 3683 627
rect -127 413 -93 447
rect -127 345 -93 379
rect -127 277 -93 311
rect -127 209 -93 243
rect -127 141 -93 175
rect -127 73 -93 107
rect 4313 413 4347 447
rect 4313 345 4347 379
rect 4313 277 4347 311
rect 4313 209 4347 243
rect 4313 141 4347 175
rect 4313 73 4347 107
rect 537 -187 571 -153
rect 605 -187 639 -153
rect 673 -187 707 -153
rect 741 -187 775 -153
rect 809 -187 843 -153
rect 1317 -187 1351 -153
rect 1385 -187 1419 -153
rect 1453 -187 1487 -153
rect 1521 -187 1555 -153
rect 1589 -187 1623 -153
rect 2597 -187 2631 -153
rect 2665 -187 2699 -153
rect 2733 -187 2767 -153
rect 2801 -187 2835 -153
rect 2869 -187 2903 -153
rect 3377 -187 3411 -153
rect 3445 -187 3479 -153
rect 3513 -187 3547 -153
rect 3581 -187 3615 -153
rect 3649 -187 3683 -153
rect -127 -447 -93 -413
rect -127 -515 -93 -481
rect -127 -583 -93 -549
rect -127 -651 -93 -617
rect -127 -719 -93 -685
rect -127 -787 -93 -753
rect 4313 -447 4347 -413
rect 4313 -515 4347 -481
rect 4313 -583 4347 -549
rect 4313 -651 4347 -617
rect 4313 -719 4347 -685
rect 4313 -787 4347 -753
rect 537 -967 571 -933
rect 605 -967 639 -933
rect 673 -967 707 -933
rect 741 -967 775 -933
rect 809 -967 843 -933
rect 1317 -967 1351 -933
rect 1385 -967 1419 -933
rect 1453 -967 1487 -933
rect 1521 -967 1555 -933
rect 1589 -967 1623 -933
rect 2597 -967 2631 -933
rect 2665 -967 2699 -933
rect 2733 -967 2767 -933
rect 2801 -967 2835 -933
rect 2869 -967 2903 -933
rect 3377 -967 3411 -933
rect 3445 -967 3479 -933
rect 3513 -967 3547 -933
rect 3581 -967 3615 -933
rect 3649 -967 3683 -933
<< locali >>
rect -140 627 4360 640
rect -140 593 529 627
rect 571 593 601 627
rect 639 593 673 627
rect 707 593 741 627
rect 779 593 809 627
rect 851 593 1309 627
rect 1351 593 1381 627
rect 1419 593 1453 627
rect 1487 593 1521 627
rect 1559 593 1589 627
rect 1631 593 2589 627
rect 2631 593 2661 627
rect 2699 593 2733 627
rect 2767 593 2801 627
rect 2839 593 2869 627
rect 2911 593 3369 627
rect 3411 593 3441 627
rect 3479 593 3513 627
rect 3547 593 3581 627
rect 3619 593 3649 627
rect 3691 593 4360 627
rect -140 580 4360 593
rect -140 447 -80 580
rect -140 413 -127 447
rect -93 413 -80 447
rect -140 379 -80 413
rect -140 345 -127 379
rect -93 345 -80 379
rect -140 311 -80 345
rect -140 277 -127 311
rect -93 277 -80 311
rect -140 243 -80 277
rect -140 209 -127 243
rect -93 209 -80 243
rect -140 175 -80 209
rect -140 141 -127 175
rect -93 141 -80 175
rect -140 107 -80 141
rect -140 73 -127 107
rect -93 73 -80 107
rect -140 -140 -80 73
rect 4300 447 4360 580
rect 4300 413 4313 447
rect 4347 413 4360 447
rect 4300 379 4360 413
rect 4300 345 4313 379
rect 4347 345 4360 379
rect 4300 311 4360 345
rect 4300 277 4313 311
rect 4347 277 4360 311
rect 4300 243 4360 277
rect 4300 209 4313 243
rect 4347 209 4360 243
rect 4300 175 4360 209
rect 4300 141 4313 175
rect 4347 141 4360 175
rect 4300 107 4360 141
rect 4300 73 4313 107
rect 4347 73 4360 107
rect 4300 -140 4360 73
rect -140 -153 4360 -140
rect -140 -187 537 -153
rect 571 -187 605 -153
rect 639 -187 673 -153
rect 707 -187 741 -153
rect 775 -187 809 -153
rect 843 -187 1317 -153
rect 1351 -187 1385 -153
rect 1419 -187 1453 -153
rect 1487 -187 1521 -153
rect 1555 -187 1589 -153
rect 1623 -187 2597 -153
rect 2631 -187 2665 -153
rect 2699 -187 2733 -153
rect 2767 -187 2801 -153
rect 2835 -187 2869 -153
rect 2903 -187 3377 -153
rect 3411 -187 3445 -153
rect 3479 -187 3513 -153
rect 3547 -187 3581 -153
rect 3615 -187 3649 -153
rect 3683 -187 4360 -153
rect -140 -200 4360 -187
rect -140 -413 -80 -200
rect -140 -447 -127 -413
rect -93 -447 -80 -413
rect -140 -481 -80 -447
rect -140 -515 -127 -481
rect -93 -515 -80 -481
rect -140 -549 -80 -515
rect -140 -583 -127 -549
rect -93 -583 -80 -549
rect -140 -617 -80 -583
rect -140 -651 -127 -617
rect -93 -651 -80 -617
rect -140 -685 -80 -651
rect -140 -719 -127 -685
rect -93 -719 -80 -685
rect -140 -753 -80 -719
rect -140 -787 -127 -753
rect -93 -787 -80 -753
rect -140 -920 -80 -787
rect 4300 -413 4360 -200
rect 4300 -447 4313 -413
rect 4347 -447 4360 -413
rect 4300 -481 4360 -447
rect 4300 -515 4313 -481
rect 4347 -515 4360 -481
rect 4300 -549 4360 -515
rect 4300 -583 4313 -549
rect 4347 -583 4360 -549
rect 4300 -617 4360 -583
rect 4300 -651 4313 -617
rect 4347 -651 4360 -617
rect 4300 -685 4360 -651
rect 4300 -719 4313 -685
rect 4347 -719 4360 -685
rect 4300 -753 4360 -719
rect 4300 -787 4313 -753
rect 4347 -787 4360 -753
rect 4300 -920 4360 -787
rect -140 -933 4360 -920
rect -140 -967 529 -933
rect 571 -967 601 -933
rect 639 -967 673 -933
rect 707 -967 741 -933
rect 779 -967 809 -933
rect 851 -967 1309 -933
rect 1351 -967 1381 -933
rect 1419 -967 1453 -933
rect 1487 -967 1521 -933
rect 1559 -967 1589 -933
rect 1631 -967 2589 -933
rect 2631 -967 2661 -933
rect 2699 -967 2733 -933
rect 2767 -967 2801 -933
rect 2839 -967 2869 -933
rect 2911 -967 3369 -933
rect 3411 -967 3441 -933
rect 3479 -967 3513 -933
rect 3547 -967 3581 -933
rect 3619 -967 3649 -933
rect 3691 -967 4360 -933
rect -140 -980 4360 -967
<< viali >>
rect 529 593 537 627
rect 537 593 563 627
rect 601 593 605 627
rect 605 593 635 627
rect 673 593 707 627
rect 745 593 775 627
rect 775 593 779 627
rect 817 593 843 627
rect 843 593 851 627
rect 1309 593 1317 627
rect 1317 593 1343 627
rect 1381 593 1385 627
rect 1385 593 1415 627
rect 1453 593 1487 627
rect 1525 593 1555 627
rect 1555 593 1559 627
rect 1597 593 1623 627
rect 1623 593 1631 627
rect 2589 593 2597 627
rect 2597 593 2623 627
rect 2661 593 2665 627
rect 2665 593 2695 627
rect 2733 593 2767 627
rect 2805 593 2835 627
rect 2835 593 2839 627
rect 2877 593 2903 627
rect 2903 593 2911 627
rect 3369 593 3377 627
rect 3377 593 3403 627
rect 3441 593 3445 627
rect 3445 593 3475 627
rect 3513 593 3547 627
rect 3585 593 3615 627
rect 3615 593 3619 627
rect 3657 593 3683 627
rect 3683 593 3691 627
rect 529 -967 537 -933
rect 537 -967 563 -933
rect 601 -967 605 -933
rect 605 -967 635 -933
rect 673 -967 707 -933
rect 745 -967 775 -933
rect 775 -967 779 -933
rect 817 -967 843 -933
rect 843 -967 851 -933
rect 1309 -967 1317 -933
rect 1317 -967 1343 -933
rect 1381 -967 1385 -933
rect 1385 -967 1415 -933
rect 1453 -967 1487 -933
rect 1525 -967 1555 -933
rect 1555 -967 1559 -933
rect 1597 -967 1623 -933
rect 1623 -967 1631 -933
rect 2589 -967 2597 -933
rect 2597 -967 2623 -933
rect 2661 -967 2665 -933
rect 2665 -967 2695 -933
rect 2733 -967 2767 -933
rect 2805 -967 2835 -933
rect 2835 -967 2839 -933
rect 2877 -967 2903 -933
rect 2903 -967 2911 -933
rect 3369 -967 3377 -933
rect 3377 -967 3403 -933
rect 3441 -967 3445 -933
rect 3445 -967 3475 -933
rect 3513 -967 3547 -933
rect 3585 -967 3615 -933
rect 3615 -967 3619 -933
rect 3657 -967 3683 -933
rect 3683 -967 3691 -933
<< metal1 >>
rect -140 627 4360 646
rect -140 593 529 627
rect 563 593 601 627
rect 635 593 673 627
rect 707 593 745 627
rect 779 593 817 627
rect 851 593 1309 627
rect 1343 593 1381 627
rect 1415 593 1453 627
rect 1487 593 1525 627
rect 1559 593 1597 627
rect 1631 593 2589 627
rect 2623 593 2661 627
rect 2695 593 2733 627
rect 2767 593 2805 627
rect 2839 593 2877 627
rect 2911 593 3369 627
rect 3403 593 3441 627
rect 3475 593 3513 627
rect 3547 593 3585 627
rect 3619 593 3657 627
rect 3691 593 4360 627
rect -140 574 4360 593
rect -140 -914 -80 574
rect 22 420 68 574
rect 538 420 584 574
rect 750 441 880 460
rect 750 389 789 441
rect 841 389 880 441
rect 1054 420 1100 574
rect 1270 441 1400 460
rect 750 370 880 389
rect 1270 389 1309 441
rect 1361 389 1400 441
rect 1570 420 1616 574
rect 2086 420 2132 574
rect 2340 448 2386 460
rect 1270 370 1400 389
rect 1316 360 1322 370
rect 1356 360 1362 370
rect 2340 150 2346 448
rect 2380 150 2386 448
rect 2598 448 2648 574
rect 240 131 370 150
rect 240 79 279 131
rect 331 79 370 131
rect 240 60 370 79
rect 1790 131 1920 150
rect 1790 79 1829 131
rect 1881 79 1920 131
rect 1790 60 1920 79
rect 2300 131 2430 150
rect 2300 79 2339 131
rect 2391 79 2430 131
rect 2300 60 2430 79
rect 2598 72 2604 448
rect 2810 441 2940 460
rect 3118 449 3164 574
rect 3330 451 3460 470
rect 2810 389 2849 441
rect 2901 389 2940 441
rect 2810 370 2940 389
rect 3330 399 3369 451
rect 3421 399 3460 451
rect 3330 380 3460 399
rect 3630 454 3680 574
rect 3888 459 3938 460
rect 3888 458 3934 459
rect 3372 370 3382 380
rect 3412 370 3422 380
rect 2856 72 2862 370
rect 2896 72 2902 370
rect 2598 60 2638 72
rect 2856 60 2902 72
rect 3372 82 3378 370
rect 3412 82 3418 370
rect 3372 70 3418 82
rect 3630 82 3636 454
rect 3670 82 3676 454
rect 3888 160 3894 458
rect 3928 160 3934 458
rect 4150 457 4196 574
rect 3630 70 3676 82
rect 3850 141 3980 160
rect 3850 89 3889 141
rect 3941 89 3980 141
rect 3850 70 3980 89
rect 280 20 330 60
rect 1830 20 1880 60
rect 2340 20 2390 60
rect 3890 20 3940 70
rect 70 -30 4140 20
rect 280 -310 330 -30
rect 1830 -310 1880 -30
rect 2340 -310 2390 -30
rect 3890 -310 3940 -30
rect 70 -360 4140 -310
rect 240 -409 370 -390
rect 240 -461 279 -409
rect 331 -461 370 -409
rect 240 -480 370 -461
rect 540 -402 586 -390
rect 282 -490 292 -480
rect 322 -490 332 -480
rect 282 -778 288 -490
rect 322 -778 328 -490
rect 21 -914 68 -789
rect 282 -790 328 -778
rect 540 -778 546 -402
rect 580 -778 586 -402
rect 798 -402 844 -390
rect 798 -700 804 -402
rect 838 -700 844 -402
rect 1310 -412 1356 -400
rect 540 -787 586 -778
rect 538 -914 586 -787
rect 760 -719 890 -700
rect 1310 -710 1316 -412
rect 1350 -710 1356 -412
rect 1568 -412 1614 -400
rect 760 -771 799 -719
rect 851 -771 890 -719
rect 760 -790 890 -771
rect 1270 -729 1400 -710
rect 1270 -781 1309 -729
rect 1361 -781 1400 -729
rect 1054 -914 1100 -789
rect 1270 -800 1400 -781
rect 1568 -788 1574 -412
rect 1608 -788 1614 -412
rect 1780 -419 1910 -400
rect 1780 -471 1819 -419
rect 1871 -471 1910 -419
rect 1780 -490 1910 -471
rect 2300 -409 2430 -390
rect 2300 -461 2339 -409
rect 2391 -461 2430 -409
rect 2300 -480 2430 -461
rect 2600 -402 2646 -390
rect 2342 -490 2352 -480
rect 2382 -490 2392 -480
rect 1568 -794 1614 -788
rect 1826 -788 1832 -490
rect 1866 -788 1872 -490
rect 1568 -914 1616 -794
rect 1826 -800 1872 -788
rect 2342 -778 2348 -490
rect 2382 -778 2388 -490
rect 2342 -790 2388 -778
rect 2600 -778 2606 -402
rect 2640 -778 2646 -402
rect 2858 -402 2904 -390
rect 2858 -700 2864 -402
rect 2898 -700 2904 -402
rect 3370 -422 3416 -410
rect 2600 -784 2646 -778
rect 2820 -719 2950 -700
rect 2820 -771 2859 -719
rect 2911 -771 2950 -719
rect 3370 -720 3376 -422
rect 3410 -720 3416 -422
rect 3628 -422 3674 -410
rect 2086 -914 2132 -794
rect 2600 -914 2648 -784
rect 2820 -790 2950 -771
rect 3330 -739 3460 -720
rect 3118 -914 3164 -778
rect 3330 -791 3369 -739
rect 3421 -791 3460 -739
rect 3330 -810 3460 -791
rect 3628 -782 3634 -422
rect 3668 -782 3674 -422
rect 3840 -429 3970 -410
rect 3840 -481 3879 -429
rect 3931 -481 3970 -429
rect 3840 -500 3970 -481
rect 3628 -914 3680 -782
rect 3886 -798 3892 -500
rect 3926 -798 3932 -500
rect 3886 -810 3932 -798
rect 4150 -914 4196 -775
rect 4300 -914 4360 574
rect -140 -933 4360 -914
rect -140 -967 529 -933
rect 563 -967 601 -933
rect 635 -967 673 -933
rect 707 -967 745 -933
rect 779 -967 817 -933
rect 851 -967 1309 -933
rect 1343 -967 1381 -933
rect 1415 -967 1453 -933
rect 1487 -967 1525 -933
rect 1559 -967 1597 -933
rect 1631 -967 2589 -933
rect 2623 -967 2661 -933
rect 2695 -967 2733 -933
rect 2767 -967 2805 -933
rect 2839 -967 2877 -933
rect 2911 -967 3369 -933
rect 3403 -967 3441 -933
rect 3475 -967 3513 -933
rect 3547 -967 3585 -933
rect 3619 -967 3657 -933
rect 3691 -967 4360 -933
rect -140 -986 4360 -967
<< via1 >>
rect 789 389 841 441
rect 1309 389 1361 441
rect 279 79 331 131
rect 1829 79 1881 131
rect 2339 79 2391 131
rect 2849 389 2901 441
rect 3369 399 3421 451
rect 3889 89 3941 141
rect 279 -461 331 -409
rect 799 -771 851 -719
rect 1309 -781 1361 -729
rect 1819 -471 1871 -419
rect 2339 -461 2391 -409
rect 2859 -771 2911 -719
rect 3369 -791 3421 -739
rect 3879 -481 3931 -429
<< metal2 >>
rect 750 451 3460 480
rect 750 443 3369 451
rect 3421 443 3460 451
rect 750 387 786 443
rect 842 441 3368 443
rect 842 389 1309 441
rect 1361 389 2849 441
rect 2901 389 3368 441
rect 842 387 3368 389
rect 3424 387 3460 443
rect 750 360 3460 387
rect 240 141 3980 170
rect 240 133 3889 141
rect 240 131 1308 133
rect 240 79 279 131
rect 331 79 1308 131
rect 240 77 1308 79
rect 1364 131 2858 133
rect 1364 79 1829 131
rect 1881 79 2339 131
rect 2391 79 2858 131
rect 1364 77 2858 79
rect 2914 89 3889 133
rect 3941 89 3980 141
rect 2914 77 3980 89
rect 240 50 3980 77
rect 250 -390 360 -380
rect 760 -390 872 -380
rect 2310 -390 2420 -380
rect 3340 -390 3452 -380
rect 240 -407 3970 -390
rect 240 -409 788 -407
rect 240 -461 279 -409
rect 331 -461 788 -409
rect 240 -463 788 -461
rect 844 -409 3368 -407
rect 844 -419 2339 -409
rect 844 -463 1819 -419
rect 240 -471 1819 -463
rect 1871 -461 2339 -419
rect 2391 -461 3368 -409
rect 1871 -463 3368 -461
rect 3424 -429 3970 -407
rect 3424 -463 3879 -429
rect 1871 -471 3879 -463
rect 240 -481 3879 -471
rect 3931 -481 3970 -429
rect 240 -490 3970 -481
rect 1790 -500 1900 -490
rect 3850 -510 3960 -490
rect 770 -710 880 -690
rect 2830 -700 2940 -690
rect 1280 -710 1392 -700
rect 2830 -710 2942 -700
rect 760 -719 3460 -710
rect 760 -771 799 -719
rect 851 -727 2859 -719
rect 2911 -727 3460 -719
rect 851 -771 1308 -727
rect 760 -783 1308 -771
rect 1364 -783 2858 -727
rect 2914 -739 3460 -727
rect 2914 -783 3369 -739
rect 760 -791 3369 -783
rect 3421 -791 3460 -739
rect 760 -810 3460 -791
rect 3340 -820 3450 -810
<< via2 >>
rect 786 441 842 443
rect 786 389 789 441
rect 789 389 841 441
rect 841 389 842 441
rect 3368 399 3369 443
rect 3369 399 3421 443
rect 3421 399 3424 443
rect 786 387 842 389
rect 3368 387 3424 399
rect 1308 77 1364 133
rect 2858 77 2914 133
rect 788 -463 844 -407
rect 3368 -463 3424 -407
rect 1308 -729 1364 -727
rect 1308 -781 1309 -729
rect 1309 -781 1361 -729
rect 1361 -781 1364 -729
rect 1308 -783 1364 -781
rect 2858 -771 2859 -727
rect 2859 -771 2911 -727
rect 2911 -771 2914 -727
rect 2858 -783 2914 -771
<< metal3 >>
rect 750 465 882 470
rect 748 443 882 465
rect 748 387 786 443
rect 842 387 882 443
rect 748 365 882 387
rect 750 -407 882 365
rect 3330 465 3460 470
rect 3330 443 3462 465
rect 3330 387 3368 443
rect 3424 387 3462 443
rect 3330 365 3462 387
rect 750 -463 788 -407
rect 844 -463 882 -407
rect 750 -490 882 -463
rect 1270 133 1402 160
rect 1270 77 1308 133
rect 1364 77 1402 133
rect 1270 -727 1402 77
rect 1270 -783 1308 -727
rect 1364 -783 1402 -727
rect 1270 -810 1402 -783
rect 2820 133 2952 155
rect 2820 77 2858 133
rect 2914 77 2952 133
rect 2820 55 2952 77
rect 2820 -705 2950 55
rect 3330 -385 3460 365
rect 3330 -407 3462 -385
rect 3330 -463 3368 -407
rect 3424 -463 3462 -407
rect 3330 -485 3462 -463
rect 2820 -727 2952 -705
rect 2820 -783 2858 -727
rect 2914 -783 2952 -727
rect 2820 -805 2952 -783
rect 2820 -810 2950 -805
rect 1270 -840 1400 -810
rect 3330 -1000 3460 -485
use sky130_fd_pr__pfet_01v8_lvt_B64SAM  sky130_fd_pr__pfet_01v8_lvt_B64SAM_0
timestamp 1663011646
transform 1 0 2109 0 1 224
box -2129 -264 2129 298
use sky130_fd_pr__pfet_01v8_lvt_MBDTEX  sky130_fd_pr__pfet_01v8_lvt_MBDTEX_0
timestamp 1663011646
transform 1 0 2109 0 1 -562
box -2129 -298 2129 264
<< end >>
