magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -226 1774 2126 1926
rect -226 -5374 -74 1774
rect 1974 -5374 2126 1774
rect -226 -5526 2126 -5374
<< psubdiff >>
rect -200 1800 2100 1900
rect -200 969 -100 1800
rect -200 935 -167 969
rect -133 935 -100 969
rect -200 901 -100 935
rect -200 867 -167 901
rect -133 867 -100 901
rect -200 833 -100 867
rect -200 799 -167 833
rect -133 799 -100 833
rect -200 765 -100 799
rect -200 731 -167 765
rect -133 731 -100 765
rect -200 -831 -100 731
rect -200 -865 -167 -831
rect -133 -865 -100 -831
rect -200 -899 -100 -865
rect -200 -933 -167 -899
rect -133 -933 -100 -899
rect -200 -967 -100 -933
rect -200 -1001 -167 -967
rect -133 -1001 -100 -967
rect -200 -1035 -100 -1001
rect -200 -1069 -167 -1035
rect -133 -1069 -100 -1035
rect -200 -2531 -100 -1069
rect -200 -2565 -167 -2531
rect -133 -2565 -100 -2531
rect -200 -2599 -100 -2565
rect -200 -2633 -167 -2599
rect -133 -2633 -100 -2599
rect -200 -2667 -100 -2633
rect -200 -2701 -167 -2667
rect -133 -2701 -100 -2667
rect -200 -2735 -100 -2701
rect -200 -2769 -167 -2735
rect -133 -2769 -100 -2735
rect -200 -4331 -100 -2769
rect -200 -4365 -167 -4331
rect -133 -4365 -100 -4331
rect -200 -4399 -100 -4365
rect -200 -4433 -167 -4399
rect -133 -4433 -100 -4399
rect -200 -4467 -100 -4433
rect -200 -4501 -167 -4467
rect -133 -4501 -100 -4467
rect -200 -4535 -100 -4501
rect -200 -4569 -167 -4535
rect -133 -4569 -100 -4535
rect -200 -5400 -100 -4569
rect 2000 969 2100 1800
rect 2000 935 2033 969
rect 2067 935 2100 969
rect 2000 901 2100 935
rect 2000 867 2033 901
rect 2067 867 2100 901
rect 2000 833 2100 867
rect 2000 799 2033 833
rect 2067 799 2100 833
rect 2000 765 2100 799
rect 2000 731 2033 765
rect 2067 731 2100 765
rect 2000 -831 2100 731
rect 2000 -865 2033 -831
rect 2067 -865 2100 -831
rect 2000 -899 2100 -865
rect 2000 -933 2033 -899
rect 2067 -933 2100 -899
rect 2000 -967 2100 -933
rect 2000 -1001 2033 -967
rect 2067 -1001 2100 -967
rect 2000 -1035 2100 -1001
rect 2000 -1069 2033 -1035
rect 2067 -1069 2100 -1035
rect 2000 -2531 2100 -1069
rect 2000 -2565 2033 -2531
rect 2067 -2565 2100 -2531
rect 2000 -2599 2100 -2565
rect 2000 -2633 2033 -2599
rect 2067 -2633 2100 -2599
rect 2000 -2667 2100 -2633
rect 2000 -2701 2033 -2667
rect 2067 -2701 2100 -2667
rect 2000 -2735 2100 -2701
rect 2000 -2769 2033 -2735
rect 2067 -2769 2100 -2735
rect 2000 -4331 2100 -2769
rect 2000 -4365 2033 -4331
rect 2067 -4365 2100 -4331
rect 2000 -4399 2100 -4365
rect 2000 -4433 2033 -4399
rect 2067 -4433 2100 -4399
rect 2000 -4467 2100 -4433
rect 2000 -4501 2033 -4467
rect 2067 -4501 2100 -4467
rect 2000 -4535 2100 -4501
rect 2000 -4569 2033 -4535
rect 2067 -4569 2100 -4535
rect 2000 -5400 2100 -4569
rect -200 -5500 2100 -5400
<< psubdiffcont >>
rect -167 935 -133 969
rect -167 867 -133 901
rect -167 799 -133 833
rect -167 731 -133 765
rect -167 -865 -133 -831
rect -167 -933 -133 -899
rect -167 -1001 -133 -967
rect -167 -1069 -133 -1035
rect -167 -2565 -133 -2531
rect -167 -2633 -133 -2599
rect -167 -2701 -133 -2667
rect -167 -2769 -133 -2735
rect -167 -4365 -133 -4331
rect -167 -4433 -133 -4399
rect -167 -4501 -133 -4467
rect -167 -4569 -133 -4535
rect 2033 935 2067 969
rect 2033 867 2067 901
rect 2033 799 2067 833
rect 2033 731 2067 765
rect 2033 -865 2067 -831
rect 2033 -933 2067 -899
rect 2033 -1001 2067 -967
rect 2033 -1069 2067 -1035
rect 2033 -2565 2067 -2531
rect 2033 -2633 2067 -2599
rect 2033 -2701 2067 -2667
rect 2033 -2769 2067 -2735
rect 2033 -4365 2067 -4331
rect 2033 -4433 2067 -4399
rect 2033 -4501 2067 -4467
rect 2033 -4569 2067 -4535
<< locali >>
rect -200 1800 2100 1900
rect -200 969 -100 1800
rect -200 935 -167 969
rect -133 935 -100 969
rect -200 901 -100 935
rect -200 867 -167 901
rect -133 867 -100 901
rect -200 833 -100 867
rect -200 799 -167 833
rect -133 799 -100 833
rect -200 765 -100 799
rect -200 731 -167 765
rect -133 731 -100 765
rect -200 -831 -100 731
rect -200 -865 -167 -831
rect -133 -865 -100 -831
rect -200 -899 -100 -865
rect -200 -933 -167 -899
rect -133 -933 -100 -899
rect -200 -967 -100 -933
rect -200 -1001 -167 -967
rect -133 -1001 -100 -967
rect -200 -1035 -100 -1001
rect -200 -1069 -167 -1035
rect -133 -1069 -100 -1035
rect -200 -2531 -100 -1069
rect -200 -2565 -167 -2531
rect -133 -2565 -100 -2531
rect -200 -2599 -100 -2565
rect -200 -2633 -167 -2599
rect -133 -2633 -100 -2599
rect -200 -2667 -100 -2633
rect -200 -2701 -167 -2667
rect -133 -2701 -100 -2667
rect -200 -2735 -100 -2701
rect -200 -2769 -167 -2735
rect -133 -2769 -100 -2735
rect -200 -4331 -100 -2769
rect -200 -4365 -167 -4331
rect -133 -4365 -100 -4331
rect -200 -4399 -100 -4365
rect -200 -4433 -167 -4399
rect -133 -4433 -100 -4399
rect -200 -4467 -100 -4433
rect -200 -4501 -167 -4467
rect -133 -4501 -100 -4467
rect -200 -4535 -100 -4501
rect -200 -4569 -167 -4535
rect -133 -4569 -100 -4535
rect -200 -5400 -100 -4569
rect 2000 969 2100 1800
rect 2000 935 2033 969
rect 2067 935 2100 969
rect 2000 901 2100 935
rect 2000 867 2033 901
rect 2067 867 2100 901
rect 2000 833 2100 867
rect 2000 799 2033 833
rect 2067 799 2100 833
rect 2000 765 2100 799
rect 2000 731 2033 765
rect 2067 731 2100 765
rect 2000 -831 2100 731
rect 2000 -865 2033 -831
rect 2067 -865 2100 -831
rect 2000 -899 2100 -865
rect 2000 -933 2033 -899
rect 2067 -933 2100 -899
rect 2000 -967 2100 -933
rect 2000 -1001 2033 -967
rect 2067 -1001 2100 -967
rect 2000 -1035 2100 -1001
rect 2000 -1069 2033 -1035
rect 2067 -1069 2100 -1035
rect 2000 -2531 2100 -1069
rect 2000 -2565 2033 -2531
rect 2067 -2565 2100 -2531
rect 2000 -2599 2100 -2565
rect 2000 -2633 2033 -2599
rect 2067 -2633 2100 -2599
rect 2000 -2667 2100 -2633
rect 2000 -2701 2033 -2667
rect 2067 -2701 2100 -2667
rect 2000 -2735 2100 -2701
rect 2000 -2769 2033 -2735
rect 2067 -2769 2100 -2735
rect 2000 -4331 2100 -2769
rect 2000 -4365 2033 -4331
rect 2067 -4365 2100 -4331
rect 2000 -4399 2100 -4365
rect 2000 -4433 2033 -4399
rect 2067 -4433 2100 -4399
rect 2000 -4467 2100 -4433
rect 2000 -4501 2033 -4467
rect 2067 -4501 2100 -4467
rect 2000 -4535 2100 -4501
rect 2000 -4569 2033 -4535
rect 2067 -4569 2100 -4535
rect 2000 -5400 2100 -4569
rect -200 -5500 2100 -5400
<< metal1 >>
rect -10 916 70 920
rect -10 864 4 916
rect 56 864 70 916
rect -10 860 70 864
rect 450 916 530 920
rect 450 864 464 916
rect 516 864 530 916
rect 450 860 530 864
rect 910 916 990 920
rect 910 864 924 916
rect 976 864 990 916
rect 910 860 990 864
rect 1370 916 1450 920
rect 1370 864 1384 916
rect 1436 864 1450 916
rect 1370 860 1450 864
rect 1830 916 1910 920
rect 1830 864 1844 916
rect 1896 864 1910 916
rect 1830 860 1910 864
rect 62 -98 1828 56
rect -10 -904 70 -900
rect -10 -956 4 -904
rect 56 -956 70 -904
rect -10 -960 70 -956
rect 450 -904 530 -900
rect 450 -956 464 -904
rect 516 -956 530 -904
rect 450 -960 530 -956
rect 910 -904 990 -900
rect 910 -956 924 -904
rect 976 -956 990 -904
rect 910 -960 990 -956
rect 1370 -904 1450 -900
rect 1370 -956 1384 -904
rect 1436 -956 1450 -904
rect 1370 -960 1450 -956
rect 1830 -904 1910 -900
rect 1830 -956 1844 -904
rect 1896 -956 1910 -904
rect 1830 -960 1910 -956
rect -10 -2584 70 -2580
rect -10 -2636 4 -2584
rect 56 -2636 70 -2584
rect -10 -2640 70 -2636
rect 450 -2584 530 -2580
rect 450 -2636 464 -2584
rect 516 -2636 530 -2584
rect 450 -2640 530 -2636
rect 910 -2584 990 -2580
rect 910 -2636 924 -2584
rect 976 -2636 990 -2584
rect 910 -2640 990 -2636
rect 1370 -2584 1450 -2580
rect 1370 -2636 1384 -2584
rect 1436 -2636 1450 -2584
rect 1370 -2640 1450 -2636
rect 1830 -2584 1910 -2580
rect 1830 -2636 1844 -2584
rect 1896 -2636 1910 -2584
rect 1830 -2640 1910 -2636
rect 62 -3610 1828 -3456
rect -10 -4404 70 -4400
rect -10 -4456 4 -4404
rect 56 -4456 70 -4404
rect -10 -4460 70 -4456
rect 450 -4404 530 -4400
rect 450 -4456 464 -4404
rect 516 -4456 530 -4404
rect 450 -4460 530 -4456
rect 910 -4404 990 -4400
rect 910 -4456 924 -4404
rect 976 -4456 990 -4404
rect 910 -4460 990 -4456
rect 1370 -4404 1450 -4400
rect 1370 -4456 1384 -4404
rect 1436 -4456 1450 -4404
rect 1370 -4460 1450 -4456
rect 1830 -4404 1910 -4400
rect 1830 -4456 1844 -4404
rect 1896 -4456 1910 -4404
rect 1830 -4460 1910 -4456
<< via1 >>
rect 4 864 56 916
rect 464 864 516 916
rect 924 864 976 916
rect 1384 864 1436 916
rect 1844 864 1896 916
rect 4 -956 56 -904
rect 464 -956 516 -904
rect 924 -956 976 -904
rect 1384 -956 1436 -904
rect 1844 -956 1896 -904
rect 4 -2636 56 -2584
rect 464 -2636 516 -2584
rect 924 -2636 976 -2584
rect 1384 -2636 1436 -2584
rect 1844 -2636 1896 -2584
rect 4 -4456 56 -4404
rect 464 -4456 516 -4404
rect 924 -4456 976 -4404
rect 1384 -4456 1436 -4404
rect 1844 -4456 1896 -4404
<< metal2 >>
rect 0 1640 1900 1700
rect 0 916 60 1640
rect 0 864 4 916
rect 56 864 60 916
rect 0 -904 60 864
rect 0 -956 4 -904
rect 56 -956 60 -904
rect 0 -970 60 -956
rect 460 916 520 930
rect 460 864 464 916
rect 516 864 520 916
rect 460 -904 520 864
rect 460 -956 464 -904
rect 516 -956 520 -904
rect 460 -1746 520 -956
rect 920 916 980 1640
rect 920 864 924 916
rect 976 864 980 916
rect 920 -904 980 864
rect 920 -956 924 -904
rect 976 -956 980 -904
rect 920 -970 980 -956
rect 1380 916 1440 930
rect 1380 864 1384 916
rect 1436 864 1440 916
rect 1380 -904 1440 864
rect 1380 -956 1384 -904
rect 1436 -956 1440 -904
rect 1380 -1746 1440 -956
rect 1840 916 1900 1640
rect 1840 864 1844 916
rect 1896 864 1900 916
rect 1840 -904 1900 864
rect 1840 -956 1844 -904
rect 1896 -956 1900 -904
rect 1840 -970 1900 -956
rect 460 -1806 1440 -1746
rect 0 -2584 60 -2570
rect 0 -2636 4 -2584
rect 56 -2636 60 -2584
rect 0 -4404 60 -2636
rect 0 -4456 4 -4404
rect 56 -4456 60 -4404
rect 0 -5180 60 -4456
rect 460 -2584 520 -1806
rect 460 -2636 464 -2584
rect 516 -2636 520 -2584
rect 460 -4404 520 -2636
rect 460 -4456 464 -4404
rect 516 -4456 520 -4404
rect 460 -4470 520 -4456
rect 920 -2584 980 -2570
rect 920 -2636 924 -2584
rect 976 -2636 980 -2584
rect 920 -4404 980 -2636
rect 920 -4456 924 -4404
rect 976 -4456 980 -4404
rect 920 -5180 980 -4456
rect 1380 -2584 1440 -1806
rect 1380 -2636 1384 -2584
rect 1436 -2636 1440 -2584
rect 1380 -4404 1440 -2636
rect 1380 -4456 1384 -4404
rect 1436 -4456 1440 -4404
rect 1380 -4470 1440 -4456
rect 1840 -2584 1900 -2570
rect 1840 -2636 1844 -2584
rect 1896 -2636 1900 -2584
rect 1840 -4404 1900 -2636
rect 1840 -4456 1844 -4404
rect 1896 -4456 1900 -4404
rect 1840 -5180 1900 -4456
rect 0 -5240 1900 -5180
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_0
timestamp 1663011646
transform 1 0 945 0 1 -899
box -971 -857 971 857
use sky130_fd_pr__nfet_01v8_lvt_64DJ5N  sky130_fd_pr__nfet_01v8_lvt_64DJ5N_1
timestamp 1663011646
transform 1 0 945 0 1 -4411
box -971 -857 971 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_0
timestamp 1663011646
transform 1 0 945 0 1 857
box -971 -857 971 857
use sky130_fd_pr__nfet_01v8_lvt_64S6GM  sky130_fd_pr__nfet_01v8_lvt_64S6GM_1
timestamp 1663011646
transform 1 0 945 0 1 -2655
box -971 -857 971 857
<< end >>
