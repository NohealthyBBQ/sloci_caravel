magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -2129 -264 2129 298
<< pmoslvt >>
rect -2035 -164 -1835 236
rect -1777 -164 -1577 236
rect -1519 -164 -1319 236
rect -1261 -164 -1061 236
rect -1003 -164 -803 236
rect -745 -164 -545 236
rect -487 -164 -287 236
rect -229 -164 -29 236
rect 29 -164 229 236
rect 287 -164 487 236
rect 545 -164 745 236
rect 803 -164 1003 236
rect 1061 -164 1261 236
rect 1319 -164 1519 236
rect 1577 -164 1777 236
rect 1835 -164 2035 236
<< pdiff >>
rect -2093 223 -2035 236
rect -2093 189 -2081 223
rect -2047 189 -2035 223
rect -2093 155 -2035 189
rect -2093 121 -2081 155
rect -2047 121 -2035 155
rect -2093 87 -2035 121
rect -2093 53 -2081 87
rect -2047 53 -2035 87
rect -2093 19 -2035 53
rect -2093 -15 -2081 19
rect -2047 -15 -2035 19
rect -2093 -49 -2035 -15
rect -2093 -83 -2081 -49
rect -2047 -83 -2035 -49
rect -2093 -117 -2035 -83
rect -2093 -151 -2081 -117
rect -2047 -151 -2035 -117
rect -2093 -164 -2035 -151
rect -1835 223 -1777 236
rect -1835 189 -1823 223
rect -1789 189 -1777 223
rect -1835 155 -1777 189
rect -1835 121 -1823 155
rect -1789 121 -1777 155
rect -1835 87 -1777 121
rect -1835 53 -1823 87
rect -1789 53 -1777 87
rect -1835 19 -1777 53
rect -1835 -15 -1823 19
rect -1789 -15 -1777 19
rect -1835 -49 -1777 -15
rect -1835 -83 -1823 -49
rect -1789 -83 -1777 -49
rect -1835 -117 -1777 -83
rect -1835 -151 -1823 -117
rect -1789 -151 -1777 -117
rect -1835 -164 -1777 -151
rect -1577 223 -1519 236
rect -1577 189 -1565 223
rect -1531 189 -1519 223
rect -1577 155 -1519 189
rect -1577 121 -1565 155
rect -1531 121 -1519 155
rect -1577 87 -1519 121
rect -1577 53 -1565 87
rect -1531 53 -1519 87
rect -1577 19 -1519 53
rect -1577 -15 -1565 19
rect -1531 -15 -1519 19
rect -1577 -49 -1519 -15
rect -1577 -83 -1565 -49
rect -1531 -83 -1519 -49
rect -1577 -117 -1519 -83
rect -1577 -151 -1565 -117
rect -1531 -151 -1519 -117
rect -1577 -164 -1519 -151
rect -1319 223 -1261 236
rect -1319 189 -1307 223
rect -1273 189 -1261 223
rect -1319 155 -1261 189
rect -1319 121 -1307 155
rect -1273 121 -1261 155
rect -1319 87 -1261 121
rect -1319 53 -1307 87
rect -1273 53 -1261 87
rect -1319 19 -1261 53
rect -1319 -15 -1307 19
rect -1273 -15 -1261 19
rect -1319 -49 -1261 -15
rect -1319 -83 -1307 -49
rect -1273 -83 -1261 -49
rect -1319 -117 -1261 -83
rect -1319 -151 -1307 -117
rect -1273 -151 -1261 -117
rect -1319 -164 -1261 -151
rect -1061 223 -1003 236
rect -1061 189 -1049 223
rect -1015 189 -1003 223
rect -1061 155 -1003 189
rect -1061 121 -1049 155
rect -1015 121 -1003 155
rect -1061 87 -1003 121
rect -1061 53 -1049 87
rect -1015 53 -1003 87
rect -1061 19 -1003 53
rect -1061 -15 -1049 19
rect -1015 -15 -1003 19
rect -1061 -49 -1003 -15
rect -1061 -83 -1049 -49
rect -1015 -83 -1003 -49
rect -1061 -117 -1003 -83
rect -1061 -151 -1049 -117
rect -1015 -151 -1003 -117
rect -1061 -164 -1003 -151
rect -803 223 -745 236
rect -803 189 -791 223
rect -757 189 -745 223
rect -803 155 -745 189
rect -803 121 -791 155
rect -757 121 -745 155
rect -803 87 -745 121
rect -803 53 -791 87
rect -757 53 -745 87
rect -803 19 -745 53
rect -803 -15 -791 19
rect -757 -15 -745 19
rect -803 -49 -745 -15
rect -803 -83 -791 -49
rect -757 -83 -745 -49
rect -803 -117 -745 -83
rect -803 -151 -791 -117
rect -757 -151 -745 -117
rect -803 -164 -745 -151
rect -545 223 -487 236
rect -545 189 -533 223
rect -499 189 -487 223
rect -545 155 -487 189
rect -545 121 -533 155
rect -499 121 -487 155
rect -545 87 -487 121
rect -545 53 -533 87
rect -499 53 -487 87
rect -545 19 -487 53
rect -545 -15 -533 19
rect -499 -15 -487 19
rect -545 -49 -487 -15
rect -545 -83 -533 -49
rect -499 -83 -487 -49
rect -545 -117 -487 -83
rect -545 -151 -533 -117
rect -499 -151 -487 -117
rect -545 -164 -487 -151
rect -287 223 -229 236
rect -287 189 -275 223
rect -241 189 -229 223
rect -287 155 -229 189
rect -287 121 -275 155
rect -241 121 -229 155
rect -287 87 -229 121
rect -287 53 -275 87
rect -241 53 -229 87
rect -287 19 -229 53
rect -287 -15 -275 19
rect -241 -15 -229 19
rect -287 -49 -229 -15
rect -287 -83 -275 -49
rect -241 -83 -229 -49
rect -287 -117 -229 -83
rect -287 -151 -275 -117
rect -241 -151 -229 -117
rect -287 -164 -229 -151
rect -29 223 29 236
rect -29 189 -17 223
rect 17 189 29 223
rect -29 155 29 189
rect -29 121 -17 155
rect 17 121 29 155
rect -29 87 29 121
rect -29 53 -17 87
rect 17 53 29 87
rect -29 19 29 53
rect -29 -15 -17 19
rect 17 -15 29 19
rect -29 -49 29 -15
rect -29 -83 -17 -49
rect 17 -83 29 -49
rect -29 -117 29 -83
rect -29 -151 -17 -117
rect 17 -151 29 -117
rect -29 -164 29 -151
rect 229 223 287 236
rect 229 189 241 223
rect 275 189 287 223
rect 229 155 287 189
rect 229 121 241 155
rect 275 121 287 155
rect 229 87 287 121
rect 229 53 241 87
rect 275 53 287 87
rect 229 19 287 53
rect 229 -15 241 19
rect 275 -15 287 19
rect 229 -49 287 -15
rect 229 -83 241 -49
rect 275 -83 287 -49
rect 229 -117 287 -83
rect 229 -151 241 -117
rect 275 -151 287 -117
rect 229 -164 287 -151
rect 487 223 545 236
rect 487 189 499 223
rect 533 189 545 223
rect 487 155 545 189
rect 487 121 499 155
rect 533 121 545 155
rect 487 87 545 121
rect 487 53 499 87
rect 533 53 545 87
rect 487 19 545 53
rect 487 -15 499 19
rect 533 -15 545 19
rect 487 -49 545 -15
rect 487 -83 499 -49
rect 533 -83 545 -49
rect 487 -117 545 -83
rect 487 -151 499 -117
rect 533 -151 545 -117
rect 487 -164 545 -151
rect 745 223 803 236
rect 745 189 757 223
rect 791 189 803 223
rect 745 155 803 189
rect 745 121 757 155
rect 791 121 803 155
rect 745 87 803 121
rect 745 53 757 87
rect 791 53 803 87
rect 745 19 803 53
rect 745 -15 757 19
rect 791 -15 803 19
rect 745 -49 803 -15
rect 745 -83 757 -49
rect 791 -83 803 -49
rect 745 -117 803 -83
rect 745 -151 757 -117
rect 791 -151 803 -117
rect 745 -164 803 -151
rect 1003 223 1061 236
rect 1003 189 1015 223
rect 1049 189 1061 223
rect 1003 155 1061 189
rect 1003 121 1015 155
rect 1049 121 1061 155
rect 1003 87 1061 121
rect 1003 53 1015 87
rect 1049 53 1061 87
rect 1003 19 1061 53
rect 1003 -15 1015 19
rect 1049 -15 1061 19
rect 1003 -49 1061 -15
rect 1003 -83 1015 -49
rect 1049 -83 1061 -49
rect 1003 -117 1061 -83
rect 1003 -151 1015 -117
rect 1049 -151 1061 -117
rect 1003 -164 1061 -151
rect 1261 223 1319 236
rect 1261 189 1273 223
rect 1307 189 1319 223
rect 1261 155 1319 189
rect 1261 121 1273 155
rect 1307 121 1319 155
rect 1261 87 1319 121
rect 1261 53 1273 87
rect 1307 53 1319 87
rect 1261 19 1319 53
rect 1261 -15 1273 19
rect 1307 -15 1319 19
rect 1261 -49 1319 -15
rect 1261 -83 1273 -49
rect 1307 -83 1319 -49
rect 1261 -117 1319 -83
rect 1261 -151 1273 -117
rect 1307 -151 1319 -117
rect 1261 -164 1319 -151
rect 1519 223 1577 236
rect 1519 189 1531 223
rect 1565 189 1577 223
rect 1519 155 1577 189
rect 1519 121 1531 155
rect 1565 121 1577 155
rect 1519 87 1577 121
rect 1519 53 1531 87
rect 1565 53 1577 87
rect 1519 19 1577 53
rect 1519 -15 1531 19
rect 1565 -15 1577 19
rect 1519 -49 1577 -15
rect 1519 -83 1531 -49
rect 1565 -83 1577 -49
rect 1519 -117 1577 -83
rect 1519 -151 1531 -117
rect 1565 -151 1577 -117
rect 1519 -164 1577 -151
rect 1777 223 1835 236
rect 1777 189 1789 223
rect 1823 189 1835 223
rect 1777 155 1835 189
rect 1777 121 1789 155
rect 1823 121 1835 155
rect 1777 87 1835 121
rect 1777 53 1789 87
rect 1823 53 1835 87
rect 1777 19 1835 53
rect 1777 -15 1789 19
rect 1823 -15 1835 19
rect 1777 -49 1835 -15
rect 1777 -83 1789 -49
rect 1823 -83 1835 -49
rect 1777 -117 1835 -83
rect 1777 -151 1789 -117
rect 1823 -151 1835 -117
rect 1777 -164 1835 -151
rect 2035 223 2093 236
rect 2035 189 2047 223
rect 2081 189 2093 223
rect 2035 155 2093 189
rect 2035 121 2047 155
rect 2081 121 2093 155
rect 2035 87 2093 121
rect 2035 53 2047 87
rect 2081 53 2093 87
rect 2035 19 2093 53
rect 2035 -15 2047 19
rect 2081 -15 2093 19
rect 2035 -49 2093 -15
rect 2035 -83 2047 -49
rect 2081 -83 2093 -49
rect 2035 -117 2093 -83
rect 2035 -151 2047 -117
rect 2081 -151 2093 -117
rect 2035 -164 2093 -151
<< pdiffc >>
rect -2081 189 -2047 223
rect -2081 121 -2047 155
rect -2081 53 -2047 87
rect -2081 -15 -2047 19
rect -2081 -83 -2047 -49
rect -2081 -151 -2047 -117
rect -1823 189 -1789 223
rect -1823 121 -1789 155
rect -1823 53 -1789 87
rect -1823 -15 -1789 19
rect -1823 -83 -1789 -49
rect -1823 -151 -1789 -117
rect -1565 189 -1531 223
rect -1565 121 -1531 155
rect -1565 53 -1531 87
rect -1565 -15 -1531 19
rect -1565 -83 -1531 -49
rect -1565 -151 -1531 -117
rect -1307 189 -1273 223
rect -1307 121 -1273 155
rect -1307 53 -1273 87
rect -1307 -15 -1273 19
rect -1307 -83 -1273 -49
rect -1307 -151 -1273 -117
rect -1049 189 -1015 223
rect -1049 121 -1015 155
rect -1049 53 -1015 87
rect -1049 -15 -1015 19
rect -1049 -83 -1015 -49
rect -1049 -151 -1015 -117
rect -791 189 -757 223
rect -791 121 -757 155
rect -791 53 -757 87
rect -791 -15 -757 19
rect -791 -83 -757 -49
rect -791 -151 -757 -117
rect -533 189 -499 223
rect -533 121 -499 155
rect -533 53 -499 87
rect -533 -15 -499 19
rect -533 -83 -499 -49
rect -533 -151 -499 -117
rect -275 189 -241 223
rect -275 121 -241 155
rect -275 53 -241 87
rect -275 -15 -241 19
rect -275 -83 -241 -49
rect -275 -151 -241 -117
rect -17 189 17 223
rect -17 121 17 155
rect -17 53 17 87
rect -17 -15 17 19
rect -17 -83 17 -49
rect -17 -151 17 -117
rect 241 189 275 223
rect 241 121 275 155
rect 241 53 275 87
rect 241 -15 275 19
rect 241 -83 275 -49
rect 241 -151 275 -117
rect 499 189 533 223
rect 499 121 533 155
rect 499 53 533 87
rect 499 -15 533 19
rect 499 -83 533 -49
rect 499 -151 533 -117
rect 757 189 791 223
rect 757 121 791 155
rect 757 53 791 87
rect 757 -15 791 19
rect 757 -83 791 -49
rect 757 -151 791 -117
rect 1015 189 1049 223
rect 1015 121 1049 155
rect 1015 53 1049 87
rect 1015 -15 1049 19
rect 1015 -83 1049 -49
rect 1015 -151 1049 -117
rect 1273 189 1307 223
rect 1273 121 1307 155
rect 1273 53 1307 87
rect 1273 -15 1307 19
rect 1273 -83 1307 -49
rect 1273 -151 1307 -117
rect 1531 189 1565 223
rect 1531 121 1565 155
rect 1531 53 1565 87
rect 1531 -15 1565 19
rect 1531 -83 1565 -49
rect 1531 -151 1565 -117
rect 1789 189 1823 223
rect 1789 121 1823 155
rect 1789 53 1823 87
rect 1789 -15 1823 19
rect 1789 -83 1823 -49
rect 1789 -151 1823 -117
rect 2047 189 2081 223
rect 2047 121 2081 155
rect 2047 53 2081 87
rect 2047 -15 2081 19
rect 2047 -83 2081 -49
rect 2047 -151 2081 -117
<< poly >>
rect -2035 236 -1835 262
rect -1777 236 -1577 262
rect -1519 236 -1319 262
rect -1261 236 -1061 262
rect -1003 236 -803 262
rect -745 236 -545 262
rect -487 236 -287 262
rect -229 236 -29 262
rect 29 236 229 262
rect 287 236 487 262
rect 545 236 745 262
rect 803 236 1003 262
rect 1061 236 1261 262
rect 1319 236 1519 262
rect 1577 236 1777 262
rect 1835 236 2035 262
rect -2035 -211 -1835 -164
rect -2035 -245 -1986 -211
rect -1952 -245 -1918 -211
rect -1884 -245 -1835 -211
rect -2035 -261 -1835 -245
rect -1777 -211 -1577 -164
rect -1777 -245 -1728 -211
rect -1694 -245 -1660 -211
rect -1626 -245 -1577 -211
rect -1777 -261 -1577 -245
rect -1519 -211 -1319 -164
rect -1519 -245 -1470 -211
rect -1436 -245 -1402 -211
rect -1368 -245 -1319 -211
rect -1519 -261 -1319 -245
rect -1261 -211 -1061 -164
rect -1261 -245 -1212 -211
rect -1178 -245 -1144 -211
rect -1110 -245 -1061 -211
rect -1261 -261 -1061 -245
rect -1003 -211 -803 -164
rect -1003 -245 -954 -211
rect -920 -245 -886 -211
rect -852 -245 -803 -211
rect -1003 -261 -803 -245
rect -745 -211 -545 -164
rect -745 -245 -696 -211
rect -662 -245 -628 -211
rect -594 -245 -545 -211
rect -745 -261 -545 -245
rect -487 -211 -287 -164
rect -487 -245 -438 -211
rect -404 -245 -370 -211
rect -336 -245 -287 -211
rect -487 -261 -287 -245
rect -229 -211 -29 -164
rect -229 -245 -180 -211
rect -146 -245 -112 -211
rect -78 -245 -29 -211
rect -229 -261 -29 -245
rect 29 -211 229 -164
rect 29 -245 78 -211
rect 112 -245 146 -211
rect 180 -245 229 -211
rect 29 -261 229 -245
rect 287 -211 487 -164
rect 287 -245 336 -211
rect 370 -245 404 -211
rect 438 -245 487 -211
rect 287 -261 487 -245
rect 545 -211 745 -164
rect 545 -245 594 -211
rect 628 -245 662 -211
rect 696 -245 745 -211
rect 545 -261 745 -245
rect 803 -211 1003 -164
rect 803 -245 852 -211
rect 886 -245 920 -211
rect 954 -245 1003 -211
rect 803 -261 1003 -245
rect 1061 -211 1261 -164
rect 1061 -245 1110 -211
rect 1144 -245 1178 -211
rect 1212 -245 1261 -211
rect 1061 -261 1261 -245
rect 1319 -211 1519 -164
rect 1319 -245 1368 -211
rect 1402 -245 1436 -211
rect 1470 -245 1519 -211
rect 1319 -261 1519 -245
rect 1577 -211 1777 -164
rect 1577 -245 1626 -211
rect 1660 -245 1694 -211
rect 1728 -245 1777 -211
rect 1577 -261 1777 -245
rect 1835 -211 2035 -164
rect 1835 -245 1884 -211
rect 1918 -245 1952 -211
rect 1986 -245 2035 -211
rect 1835 -261 2035 -245
<< polycont >>
rect -1986 -245 -1952 -211
rect -1918 -245 -1884 -211
rect -1728 -245 -1694 -211
rect -1660 -245 -1626 -211
rect -1470 -245 -1436 -211
rect -1402 -245 -1368 -211
rect -1212 -245 -1178 -211
rect -1144 -245 -1110 -211
rect -954 -245 -920 -211
rect -886 -245 -852 -211
rect -696 -245 -662 -211
rect -628 -245 -594 -211
rect -438 -245 -404 -211
rect -370 -245 -336 -211
rect -180 -245 -146 -211
rect -112 -245 -78 -211
rect 78 -245 112 -211
rect 146 -245 180 -211
rect 336 -245 370 -211
rect 404 -245 438 -211
rect 594 -245 628 -211
rect 662 -245 696 -211
rect 852 -245 886 -211
rect 920 -245 954 -211
rect 1110 -245 1144 -211
rect 1178 -245 1212 -211
rect 1368 -245 1402 -211
rect 1436 -245 1470 -211
rect 1626 -245 1660 -211
rect 1694 -245 1728 -211
rect 1884 -245 1918 -211
rect 1952 -245 1986 -211
<< locali >>
rect -2081 223 -2047 240
rect -2081 155 -2047 163
rect -2081 87 -2047 91
rect -2081 -19 -2047 -15
rect -2081 -91 -2047 -83
rect -2081 -168 -2047 -151
rect -1823 223 -1789 240
rect -1823 155 -1789 163
rect -1823 87 -1789 91
rect -1823 -19 -1789 -15
rect -1823 -91 -1789 -83
rect -1823 -168 -1789 -151
rect -1565 223 -1531 240
rect -1565 155 -1531 163
rect -1565 87 -1531 91
rect -1565 -19 -1531 -15
rect -1565 -91 -1531 -83
rect -1565 -168 -1531 -151
rect -1307 223 -1273 240
rect -1307 155 -1273 163
rect -1307 87 -1273 91
rect -1307 -19 -1273 -15
rect -1307 -91 -1273 -83
rect -1307 -168 -1273 -151
rect -1049 223 -1015 240
rect -1049 155 -1015 163
rect -1049 87 -1015 91
rect -1049 -19 -1015 -15
rect -1049 -91 -1015 -83
rect -1049 -168 -1015 -151
rect -791 223 -757 240
rect -791 155 -757 163
rect -791 87 -757 91
rect -791 -19 -757 -15
rect -791 -91 -757 -83
rect -791 -168 -757 -151
rect -533 223 -499 240
rect -533 155 -499 163
rect -533 87 -499 91
rect -533 -19 -499 -15
rect -533 -91 -499 -83
rect -533 -168 -499 -151
rect -275 223 -241 240
rect -275 155 -241 163
rect -275 87 -241 91
rect -275 -19 -241 -15
rect -275 -91 -241 -83
rect -275 -168 -241 -151
rect -17 223 17 240
rect -17 155 17 163
rect -17 87 17 91
rect -17 -19 17 -15
rect -17 -91 17 -83
rect -17 -168 17 -151
rect 241 223 275 240
rect 241 155 275 163
rect 241 87 275 91
rect 241 -19 275 -15
rect 241 -91 275 -83
rect 241 -168 275 -151
rect 499 223 533 240
rect 499 155 533 163
rect 499 87 533 91
rect 499 -19 533 -15
rect 499 -91 533 -83
rect 499 -168 533 -151
rect 757 223 791 240
rect 757 155 791 163
rect 757 87 791 91
rect 757 -19 791 -15
rect 757 -91 791 -83
rect 757 -168 791 -151
rect 1015 223 1049 240
rect 1015 155 1049 163
rect 1015 87 1049 91
rect 1015 -19 1049 -15
rect 1015 -91 1049 -83
rect 1015 -168 1049 -151
rect 1273 223 1307 240
rect 1273 155 1307 163
rect 1273 87 1307 91
rect 1273 -19 1307 -15
rect 1273 -91 1307 -83
rect 1273 -168 1307 -151
rect 1531 223 1565 240
rect 1531 155 1565 163
rect 1531 87 1565 91
rect 1531 -19 1565 -15
rect 1531 -91 1565 -83
rect 1531 -168 1565 -151
rect 1789 223 1823 240
rect 1789 155 1823 163
rect 1789 87 1823 91
rect 1789 -19 1823 -15
rect 1789 -91 1823 -83
rect 1789 -168 1823 -151
rect 2047 223 2081 240
rect 2047 155 2081 163
rect 2047 87 2081 91
rect 2047 -19 2081 -15
rect 2047 -91 2081 -83
rect 2047 -168 2081 -151
rect -2035 -245 -1988 -211
rect -1952 -245 -1918 -211
rect -1882 -245 -1835 -211
rect -1777 -245 -1730 -211
rect -1694 -245 -1660 -211
rect -1624 -245 -1577 -211
rect -1519 -245 -1472 -211
rect -1436 -245 -1402 -211
rect -1366 -245 -1319 -211
rect -1261 -245 -1214 -211
rect -1178 -245 -1144 -211
rect -1108 -245 -1061 -211
rect -1003 -245 -956 -211
rect -920 -245 -886 -211
rect -850 -245 -803 -211
rect -745 -245 -698 -211
rect -662 -245 -628 -211
rect -592 -245 -545 -211
rect -487 -245 -440 -211
rect -404 -245 -370 -211
rect -334 -245 -287 -211
rect -229 -245 -182 -211
rect -146 -245 -112 -211
rect -76 -245 -29 -211
rect 29 -245 76 -211
rect 112 -245 146 -211
rect 182 -245 229 -211
rect 287 -245 334 -211
rect 370 -245 404 -211
rect 440 -245 487 -211
rect 545 -245 592 -211
rect 628 -245 662 -211
rect 698 -245 745 -211
rect 803 -245 850 -211
rect 886 -245 920 -211
rect 956 -245 1003 -211
rect 1061 -245 1108 -211
rect 1144 -245 1178 -211
rect 1214 -245 1261 -211
rect 1319 -245 1366 -211
rect 1402 -245 1436 -211
rect 1472 -245 1519 -211
rect 1577 -245 1624 -211
rect 1660 -245 1694 -211
rect 1730 -245 1777 -211
rect 1835 -245 1882 -211
rect 1918 -245 1952 -211
rect 1988 -245 2035 -211
<< viali >>
rect -2081 189 -2047 197
rect -2081 163 -2047 189
rect -2081 121 -2047 125
rect -2081 91 -2047 121
rect -2081 19 -2047 53
rect -2081 -49 -2047 -19
rect -2081 -53 -2047 -49
rect -2081 -117 -2047 -91
rect -2081 -125 -2047 -117
rect -1823 189 -1789 197
rect -1823 163 -1789 189
rect -1823 121 -1789 125
rect -1823 91 -1789 121
rect -1823 19 -1789 53
rect -1823 -49 -1789 -19
rect -1823 -53 -1789 -49
rect -1823 -117 -1789 -91
rect -1823 -125 -1789 -117
rect -1565 189 -1531 197
rect -1565 163 -1531 189
rect -1565 121 -1531 125
rect -1565 91 -1531 121
rect -1565 19 -1531 53
rect -1565 -49 -1531 -19
rect -1565 -53 -1531 -49
rect -1565 -117 -1531 -91
rect -1565 -125 -1531 -117
rect -1307 189 -1273 197
rect -1307 163 -1273 189
rect -1307 121 -1273 125
rect -1307 91 -1273 121
rect -1307 19 -1273 53
rect -1307 -49 -1273 -19
rect -1307 -53 -1273 -49
rect -1307 -117 -1273 -91
rect -1307 -125 -1273 -117
rect -1049 189 -1015 197
rect -1049 163 -1015 189
rect -1049 121 -1015 125
rect -1049 91 -1015 121
rect -1049 19 -1015 53
rect -1049 -49 -1015 -19
rect -1049 -53 -1015 -49
rect -1049 -117 -1015 -91
rect -1049 -125 -1015 -117
rect -791 189 -757 197
rect -791 163 -757 189
rect -791 121 -757 125
rect -791 91 -757 121
rect -791 19 -757 53
rect -791 -49 -757 -19
rect -791 -53 -757 -49
rect -791 -117 -757 -91
rect -791 -125 -757 -117
rect -533 189 -499 197
rect -533 163 -499 189
rect -533 121 -499 125
rect -533 91 -499 121
rect -533 19 -499 53
rect -533 -49 -499 -19
rect -533 -53 -499 -49
rect -533 -117 -499 -91
rect -533 -125 -499 -117
rect -275 189 -241 197
rect -275 163 -241 189
rect -275 121 -241 125
rect -275 91 -241 121
rect -275 19 -241 53
rect -275 -49 -241 -19
rect -275 -53 -241 -49
rect -275 -117 -241 -91
rect -275 -125 -241 -117
rect -17 189 17 197
rect -17 163 17 189
rect -17 121 17 125
rect -17 91 17 121
rect -17 19 17 53
rect -17 -49 17 -19
rect -17 -53 17 -49
rect -17 -117 17 -91
rect -17 -125 17 -117
rect 241 189 275 197
rect 241 163 275 189
rect 241 121 275 125
rect 241 91 275 121
rect 241 19 275 53
rect 241 -49 275 -19
rect 241 -53 275 -49
rect 241 -117 275 -91
rect 241 -125 275 -117
rect 499 189 533 197
rect 499 163 533 189
rect 499 121 533 125
rect 499 91 533 121
rect 499 19 533 53
rect 499 -49 533 -19
rect 499 -53 533 -49
rect 499 -117 533 -91
rect 499 -125 533 -117
rect 757 189 791 197
rect 757 163 791 189
rect 757 121 791 125
rect 757 91 791 121
rect 757 19 791 53
rect 757 -49 791 -19
rect 757 -53 791 -49
rect 757 -117 791 -91
rect 757 -125 791 -117
rect 1015 189 1049 197
rect 1015 163 1049 189
rect 1015 121 1049 125
rect 1015 91 1049 121
rect 1015 19 1049 53
rect 1015 -49 1049 -19
rect 1015 -53 1049 -49
rect 1015 -117 1049 -91
rect 1015 -125 1049 -117
rect 1273 189 1307 197
rect 1273 163 1307 189
rect 1273 121 1307 125
rect 1273 91 1307 121
rect 1273 19 1307 53
rect 1273 -49 1307 -19
rect 1273 -53 1307 -49
rect 1273 -117 1307 -91
rect 1273 -125 1307 -117
rect 1531 189 1565 197
rect 1531 163 1565 189
rect 1531 121 1565 125
rect 1531 91 1565 121
rect 1531 19 1565 53
rect 1531 -49 1565 -19
rect 1531 -53 1565 -49
rect 1531 -117 1565 -91
rect 1531 -125 1565 -117
rect 1789 189 1823 197
rect 1789 163 1823 189
rect 1789 121 1823 125
rect 1789 91 1823 121
rect 1789 19 1823 53
rect 1789 -49 1823 -19
rect 1789 -53 1823 -49
rect 1789 -117 1823 -91
rect 1789 -125 1823 -117
rect 2047 189 2081 197
rect 2047 163 2081 189
rect 2047 121 2081 125
rect 2047 91 2081 121
rect 2047 19 2081 53
rect 2047 -49 2081 -19
rect 2047 -53 2081 -49
rect 2047 -117 2081 -91
rect 2047 -125 2081 -117
rect -1988 -245 -1986 -211
rect -1986 -245 -1954 -211
rect -1916 -245 -1884 -211
rect -1884 -245 -1882 -211
rect -1730 -245 -1728 -211
rect -1728 -245 -1696 -211
rect -1658 -245 -1626 -211
rect -1626 -245 -1624 -211
rect -1472 -245 -1470 -211
rect -1470 -245 -1438 -211
rect -1400 -245 -1368 -211
rect -1368 -245 -1366 -211
rect -1214 -245 -1212 -211
rect -1212 -245 -1180 -211
rect -1142 -245 -1110 -211
rect -1110 -245 -1108 -211
rect -956 -245 -954 -211
rect -954 -245 -922 -211
rect -884 -245 -852 -211
rect -852 -245 -850 -211
rect -698 -245 -696 -211
rect -696 -245 -664 -211
rect -626 -245 -594 -211
rect -594 -245 -592 -211
rect -440 -245 -438 -211
rect -438 -245 -406 -211
rect -368 -245 -336 -211
rect -336 -245 -334 -211
rect -182 -245 -180 -211
rect -180 -245 -148 -211
rect -110 -245 -78 -211
rect -78 -245 -76 -211
rect 76 -245 78 -211
rect 78 -245 110 -211
rect 148 -245 180 -211
rect 180 -245 182 -211
rect 334 -245 336 -211
rect 336 -245 368 -211
rect 406 -245 438 -211
rect 438 -245 440 -211
rect 592 -245 594 -211
rect 594 -245 626 -211
rect 664 -245 696 -211
rect 696 -245 698 -211
rect 850 -245 852 -211
rect 852 -245 884 -211
rect 922 -245 954 -211
rect 954 -245 956 -211
rect 1108 -245 1110 -211
rect 1110 -245 1142 -211
rect 1180 -245 1212 -211
rect 1212 -245 1214 -211
rect 1366 -245 1368 -211
rect 1368 -245 1400 -211
rect 1438 -245 1470 -211
rect 1470 -245 1472 -211
rect 1624 -245 1626 -211
rect 1626 -245 1658 -211
rect 1696 -245 1728 -211
rect 1728 -245 1730 -211
rect 1882 -245 1884 -211
rect 1884 -245 1916 -211
rect 1954 -245 1986 -211
rect 1986 -245 1988 -211
<< metal1 >>
rect -2087 197 -2041 236
rect -2087 163 -2081 197
rect -2047 163 -2041 197
rect -2087 125 -2041 163
rect -2087 91 -2081 125
rect -2047 91 -2041 125
rect -2087 53 -2041 91
rect -2087 19 -2081 53
rect -2047 19 -2041 53
rect -2087 -19 -2041 19
rect -2087 -53 -2081 -19
rect -2047 -53 -2041 -19
rect -2087 -91 -2041 -53
rect -2087 -125 -2081 -91
rect -2047 -125 -2041 -91
rect -2087 -164 -2041 -125
rect -1829 197 -1783 236
rect -1829 163 -1823 197
rect -1789 163 -1783 197
rect -1829 125 -1783 163
rect -1829 91 -1823 125
rect -1789 91 -1783 125
rect -1829 53 -1783 91
rect -1829 19 -1823 53
rect -1789 19 -1783 53
rect -1829 -19 -1783 19
rect -1829 -53 -1823 -19
rect -1789 -53 -1783 -19
rect -1829 -91 -1783 -53
rect -1829 -125 -1823 -91
rect -1789 -125 -1783 -91
rect -1829 -164 -1783 -125
rect -1571 197 -1525 236
rect -1571 163 -1565 197
rect -1531 163 -1525 197
rect -1571 125 -1525 163
rect -1571 91 -1565 125
rect -1531 91 -1525 125
rect -1571 53 -1525 91
rect -1571 19 -1565 53
rect -1531 19 -1525 53
rect -1571 -19 -1525 19
rect -1571 -53 -1565 -19
rect -1531 -53 -1525 -19
rect -1571 -91 -1525 -53
rect -1571 -125 -1565 -91
rect -1531 -125 -1525 -91
rect -1571 -164 -1525 -125
rect -1313 197 -1267 236
rect -1313 163 -1307 197
rect -1273 163 -1267 197
rect -1313 125 -1267 163
rect -1313 91 -1307 125
rect -1273 91 -1267 125
rect -1313 53 -1267 91
rect -1313 19 -1307 53
rect -1273 19 -1267 53
rect -1313 -19 -1267 19
rect -1313 -53 -1307 -19
rect -1273 -53 -1267 -19
rect -1313 -91 -1267 -53
rect -1313 -125 -1307 -91
rect -1273 -125 -1267 -91
rect -1313 -164 -1267 -125
rect -1055 197 -1009 236
rect -1055 163 -1049 197
rect -1015 163 -1009 197
rect -1055 125 -1009 163
rect -1055 91 -1049 125
rect -1015 91 -1009 125
rect -1055 53 -1009 91
rect -1055 19 -1049 53
rect -1015 19 -1009 53
rect -1055 -19 -1009 19
rect -1055 -53 -1049 -19
rect -1015 -53 -1009 -19
rect -1055 -91 -1009 -53
rect -1055 -125 -1049 -91
rect -1015 -125 -1009 -91
rect -1055 -164 -1009 -125
rect -797 197 -751 236
rect -797 163 -791 197
rect -757 163 -751 197
rect -797 125 -751 163
rect -797 91 -791 125
rect -757 91 -751 125
rect -797 53 -751 91
rect -797 19 -791 53
rect -757 19 -751 53
rect -797 -19 -751 19
rect -797 -53 -791 -19
rect -757 -53 -751 -19
rect -797 -91 -751 -53
rect -797 -125 -791 -91
rect -757 -125 -751 -91
rect -797 -164 -751 -125
rect -539 197 -493 236
rect -539 163 -533 197
rect -499 163 -493 197
rect -539 125 -493 163
rect -539 91 -533 125
rect -499 91 -493 125
rect -539 53 -493 91
rect -539 19 -533 53
rect -499 19 -493 53
rect -539 -19 -493 19
rect -539 -53 -533 -19
rect -499 -53 -493 -19
rect -539 -91 -493 -53
rect -539 -125 -533 -91
rect -499 -125 -493 -91
rect -539 -164 -493 -125
rect -281 197 -235 236
rect -281 163 -275 197
rect -241 163 -235 197
rect -281 125 -235 163
rect -281 91 -275 125
rect -241 91 -235 125
rect -281 53 -235 91
rect -281 19 -275 53
rect -241 19 -235 53
rect -281 -19 -235 19
rect -281 -53 -275 -19
rect -241 -53 -235 -19
rect -281 -91 -235 -53
rect -281 -125 -275 -91
rect -241 -125 -235 -91
rect -281 -164 -235 -125
rect -23 197 23 236
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -164 23 -125
rect 235 197 281 236
rect 235 163 241 197
rect 275 163 281 197
rect 235 125 281 163
rect 235 91 241 125
rect 275 91 281 125
rect 235 53 281 91
rect 235 19 241 53
rect 275 19 281 53
rect 235 -19 281 19
rect 235 -53 241 -19
rect 275 -53 281 -19
rect 235 -91 281 -53
rect 235 -125 241 -91
rect 275 -125 281 -91
rect 235 -164 281 -125
rect 493 197 539 236
rect 493 163 499 197
rect 533 163 539 197
rect 493 125 539 163
rect 493 91 499 125
rect 533 91 539 125
rect 493 53 539 91
rect 493 19 499 53
rect 533 19 539 53
rect 493 -19 539 19
rect 493 -53 499 -19
rect 533 -53 539 -19
rect 493 -91 539 -53
rect 493 -125 499 -91
rect 533 -125 539 -91
rect 493 -164 539 -125
rect 751 197 797 236
rect 751 163 757 197
rect 791 163 797 197
rect 751 125 797 163
rect 751 91 757 125
rect 791 91 797 125
rect 751 53 797 91
rect 751 19 757 53
rect 791 19 797 53
rect 751 -19 797 19
rect 751 -53 757 -19
rect 791 -53 797 -19
rect 751 -91 797 -53
rect 751 -125 757 -91
rect 791 -125 797 -91
rect 751 -164 797 -125
rect 1009 197 1055 236
rect 1009 163 1015 197
rect 1049 163 1055 197
rect 1009 125 1055 163
rect 1009 91 1015 125
rect 1049 91 1055 125
rect 1009 53 1055 91
rect 1009 19 1015 53
rect 1049 19 1055 53
rect 1009 -19 1055 19
rect 1009 -53 1015 -19
rect 1049 -53 1055 -19
rect 1009 -91 1055 -53
rect 1009 -125 1015 -91
rect 1049 -125 1055 -91
rect 1009 -164 1055 -125
rect 1267 197 1313 236
rect 1267 163 1273 197
rect 1307 163 1313 197
rect 1267 125 1313 163
rect 1267 91 1273 125
rect 1307 91 1313 125
rect 1267 53 1313 91
rect 1267 19 1273 53
rect 1307 19 1313 53
rect 1267 -19 1313 19
rect 1267 -53 1273 -19
rect 1307 -53 1313 -19
rect 1267 -91 1313 -53
rect 1267 -125 1273 -91
rect 1307 -125 1313 -91
rect 1267 -164 1313 -125
rect 1525 197 1571 236
rect 1525 163 1531 197
rect 1565 163 1571 197
rect 1525 125 1571 163
rect 1525 91 1531 125
rect 1565 91 1571 125
rect 1525 53 1571 91
rect 1525 19 1531 53
rect 1565 19 1571 53
rect 1525 -19 1571 19
rect 1525 -53 1531 -19
rect 1565 -53 1571 -19
rect 1525 -91 1571 -53
rect 1525 -125 1531 -91
rect 1565 -125 1571 -91
rect 1525 -164 1571 -125
rect 1783 197 1829 236
rect 1783 163 1789 197
rect 1823 163 1829 197
rect 1783 125 1829 163
rect 1783 91 1789 125
rect 1823 91 1829 125
rect 1783 53 1829 91
rect 1783 19 1789 53
rect 1823 19 1829 53
rect 1783 -19 1829 19
rect 1783 -53 1789 -19
rect 1823 -53 1829 -19
rect 1783 -91 1829 -53
rect 1783 -125 1789 -91
rect 1823 -125 1829 -91
rect 1783 -164 1829 -125
rect 2041 197 2087 236
rect 2041 163 2047 197
rect 2081 163 2087 197
rect 2041 125 2087 163
rect 2041 91 2047 125
rect 2081 91 2087 125
rect 2041 53 2087 91
rect 2041 19 2047 53
rect 2081 19 2087 53
rect 2041 -19 2087 19
rect 2041 -53 2047 -19
rect 2081 -53 2087 -19
rect 2041 -91 2087 -53
rect 2041 -125 2047 -91
rect 2081 -125 2087 -91
rect 2041 -164 2087 -125
rect -2031 -211 -1839 -205
rect -2031 -245 -1988 -211
rect -1954 -245 -1916 -211
rect -1882 -245 -1839 -211
rect -2031 -251 -1839 -245
rect -1773 -211 -1581 -205
rect -1773 -245 -1730 -211
rect -1696 -245 -1658 -211
rect -1624 -245 -1581 -211
rect -1773 -251 -1581 -245
rect -1515 -211 -1323 -205
rect -1515 -245 -1472 -211
rect -1438 -245 -1400 -211
rect -1366 -245 -1323 -211
rect -1515 -251 -1323 -245
rect -1257 -211 -1065 -205
rect -1257 -245 -1214 -211
rect -1180 -245 -1142 -211
rect -1108 -245 -1065 -211
rect -1257 -251 -1065 -245
rect -999 -211 -807 -205
rect -999 -245 -956 -211
rect -922 -245 -884 -211
rect -850 -245 -807 -211
rect -999 -251 -807 -245
rect -741 -211 -549 -205
rect -741 -245 -698 -211
rect -664 -245 -626 -211
rect -592 -245 -549 -211
rect -741 -251 -549 -245
rect -483 -211 -291 -205
rect -483 -245 -440 -211
rect -406 -245 -368 -211
rect -334 -245 -291 -211
rect -483 -251 -291 -245
rect -225 -211 -33 -205
rect -225 -245 -182 -211
rect -148 -245 -110 -211
rect -76 -245 -33 -211
rect -225 -251 -33 -245
rect 33 -211 225 -205
rect 33 -245 76 -211
rect 110 -245 148 -211
rect 182 -245 225 -211
rect 33 -251 225 -245
rect 291 -211 483 -205
rect 291 -245 334 -211
rect 368 -245 406 -211
rect 440 -245 483 -211
rect 291 -251 483 -245
rect 549 -211 741 -205
rect 549 -245 592 -211
rect 626 -245 664 -211
rect 698 -245 741 -211
rect 549 -251 741 -245
rect 807 -211 999 -205
rect 807 -245 850 -211
rect 884 -245 922 -211
rect 956 -245 999 -211
rect 807 -251 999 -245
rect 1065 -211 1257 -205
rect 1065 -245 1108 -211
rect 1142 -245 1180 -211
rect 1214 -245 1257 -211
rect 1065 -251 1257 -245
rect 1323 -211 1515 -205
rect 1323 -245 1366 -211
rect 1400 -245 1438 -211
rect 1472 -245 1515 -211
rect 1323 -251 1515 -245
rect 1581 -211 1773 -205
rect 1581 -245 1624 -211
rect 1658 -245 1696 -211
rect 1730 -245 1773 -211
rect 1581 -251 1773 -245
rect 1839 -211 2031 -205
rect 1839 -245 1882 -211
rect 1916 -245 1954 -211
rect 1988 -245 2031 -211
rect 1839 -251 2031 -245
<< end >>
