magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -927 181 -865 187
rect -799 181 -737 187
rect -671 181 -609 187
rect -543 181 -481 187
rect -415 181 -353 187
rect -287 181 -225 187
rect -159 181 -97 187
rect -31 181 31 187
rect 97 181 159 187
rect 225 181 287 187
rect 353 181 415 187
rect 481 181 543 187
rect 609 181 671 187
rect 737 181 799 187
rect 865 181 927 187
rect -927 147 -913 181
rect -799 147 -785 181
rect -671 147 -657 181
rect -543 147 -529 181
rect -415 147 -401 181
rect -287 147 -273 181
rect -159 147 -145 181
rect -31 147 -17 181
rect 97 147 111 181
rect 225 147 239 181
rect 353 147 367 181
rect 481 147 495 181
rect 609 147 623 181
rect 737 147 751 181
rect 865 147 879 181
rect -927 141 -865 147
rect -799 141 -737 147
rect -671 141 -609 147
rect -543 141 -481 147
rect -415 141 -353 147
rect -287 141 -225 147
rect -159 141 -97 147
rect -31 141 31 147
rect 97 141 159 147
rect 225 141 287 147
rect 353 141 415 147
rect 481 141 543 147
rect 609 141 671 147
rect 737 141 799 147
rect 865 141 927 147
rect -927 -147 -865 -141
rect -799 -147 -737 -141
rect -671 -147 -609 -141
rect -543 -147 -481 -141
rect -415 -147 -353 -141
rect -287 -147 -225 -141
rect -159 -147 -97 -141
rect -31 -147 31 -141
rect 97 -147 159 -141
rect 225 -147 287 -141
rect 353 -147 415 -141
rect 481 -147 543 -141
rect 609 -147 671 -141
rect 737 -147 799 -141
rect 865 -147 927 -141
rect -927 -181 -913 -147
rect -799 -181 -785 -147
rect -671 -181 -657 -147
rect -543 -181 -529 -147
rect -415 -181 -401 -147
rect -287 -181 -273 -147
rect -159 -181 -145 -147
rect -31 -181 -17 -147
rect 97 -181 111 -147
rect 225 -181 239 -147
rect 353 -181 367 -147
rect 481 -181 495 -147
rect 609 -181 623 -147
rect 737 -181 751 -147
rect 865 -181 879 -147
rect -927 -187 -865 -181
rect -799 -187 -737 -181
rect -671 -187 -609 -181
rect -543 -187 -481 -181
rect -415 -187 -353 -181
rect -287 -187 -225 -181
rect -159 -187 -97 -181
rect -31 -187 31 -181
rect 97 -187 159 -181
rect 225 -187 287 -181
rect 353 -187 415 -181
rect 481 -187 543 -181
rect 609 -187 671 -181
rect 737 -187 799 -181
rect 865 -187 927 -181
<< nwell >>
rect -1127 -319 1127 319
<< pmoslvt >>
rect -931 -100 -861 100
rect -803 -100 -733 100
rect -675 -100 -605 100
rect -547 -100 -477 100
rect -419 -100 -349 100
rect -291 -100 -221 100
rect -163 -100 -93 100
rect -35 -100 35 100
rect 93 -100 163 100
rect 221 -100 291 100
rect 349 -100 419 100
rect 477 -100 547 100
rect 605 -100 675 100
rect 733 -100 803 100
rect 861 -100 931 100
<< pdiff >>
rect -989 85 -931 100
rect -989 51 -977 85
rect -943 51 -931 85
rect -989 17 -931 51
rect -989 -17 -977 17
rect -943 -17 -931 17
rect -989 -51 -931 -17
rect -989 -85 -977 -51
rect -943 -85 -931 -51
rect -989 -100 -931 -85
rect -861 85 -803 100
rect -861 51 -849 85
rect -815 51 -803 85
rect -861 17 -803 51
rect -861 -17 -849 17
rect -815 -17 -803 17
rect -861 -51 -803 -17
rect -861 -85 -849 -51
rect -815 -85 -803 -51
rect -861 -100 -803 -85
rect -733 85 -675 100
rect -733 51 -721 85
rect -687 51 -675 85
rect -733 17 -675 51
rect -733 -17 -721 17
rect -687 -17 -675 17
rect -733 -51 -675 -17
rect -733 -85 -721 -51
rect -687 -85 -675 -51
rect -733 -100 -675 -85
rect -605 85 -547 100
rect -605 51 -593 85
rect -559 51 -547 85
rect -605 17 -547 51
rect -605 -17 -593 17
rect -559 -17 -547 17
rect -605 -51 -547 -17
rect -605 -85 -593 -51
rect -559 -85 -547 -51
rect -605 -100 -547 -85
rect -477 85 -419 100
rect -477 51 -465 85
rect -431 51 -419 85
rect -477 17 -419 51
rect -477 -17 -465 17
rect -431 -17 -419 17
rect -477 -51 -419 -17
rect -477 -85 -465 -51
rect -431 -85 -419 -51
rect -477 -100 -419 -85
rect -349 85 -291 100
rect -349 51 -337 85
rect -303 51 -291 85
rect -349 17 -291 51
rect -349 -17 -337 17
rect -303 -17 -291 17
rect -349 -51 -291 -17
rect -349 -85 -337 -51
rect -303 -85 -291 -51
rect -349 -100 -291 -85
rect -221 85 -163 100
rect -221 51 -209 85
rect -175 51 -163 85
rect -221 17 -163 51
rect -221 -17 -209 17
rect -175 -17 -163 17
rect -221 -51 -163 -17
rect -221 -85 -209 -51
rect -175 -85 -163 -51
rect -221 -100 -163 -85
rect -93 85 -35 100
rect -93 51 -81 85
rect -47 51 -35 85
rect -93 17 -35 51
rect -93 -17 -81 17
rect -47 -17 -35 17
rect -93 -51 -35 -17
rect -93 -85 -81 -51
rect -47 -85 -35 -51
rect -93 -100 -35 -85
rect 35 85 93 100
rect 35 51 47 85
rect 81 51 93 85
rect 35 17 93 51
rect 35 -17 47 17
rect 81 -17 93 17
rect 35 -51 93 -17
rect 35 -85 47 -51
rect 81 -85 93 -51
rect 35 -100 93 -85
rect 163 85 221 100
rect 163 51 175 85
rect 209 51 221 85
rect 163 17 221 51
rect 163 -17 175 17
rect 209 -17 221 17
rect 163 -51 221 -17
rect 163 -85 175 -51
rect 209 -85 221 -51
rect 163 -100 221 -85
rect 291 85 349 100
rect 291 51 303 85
rect 337 51 349 85
rect 291 17 349 51
rect 291 -17 303 17
rect 337 -17 349 17
rect 291 -51 349 -17
rect 291 -85 303 -51
rect 337 -85 349 -51
rect 291 -100 349 -85
rect 419 85 477 100
rect 419 51 431 85
rect 465 51 477 85
rect 419 17 477 51
rect 419 -17 431 17
rect 465 -17 477 17
rect 419 -51 477 -17
rect 419 -85 431 -51
rect 465 -85 477 -51
rect 419 -100 477 -85
rect 547 85 605 100
rect 547 51 559 85
rect 593 51 605 85
rect 547 17 605 51
rect 547 -17 559 17
rect 593 -17 605 17
rect 547 -51 605 -17
rect 547 -85 559 -51
rect 593 -85 605 -51
rect 547 -100 605 -85
rect 675 85 733 100
rect 675 51 687 85
rect 721 51 733 85
rect 675 17 733 51
rect 675 -17 687 17
rect 721 -17 733 17
rect 675 -51 733 -17
rect 675 -85 687 -51
rect 721 -85 733 -51
rect 675 -100 733 -85
rect 803 85 861 100
rect 803 51 815 85
rect 849 51 861 85
rect 803 17 861 51
rect 803 -17 815 17
rect 849 -17 861 17
rect 803 -51 861 -17
rect 803 -85 815 -51
rect 849 -85 861 -51
rect 803 -100 861 -85
rect 931 85 989 100
rect 931 51 943 85
rect 977 51 989 85
rect 931 17 989 51
rect 931 -17 943 17
rect 977 -17 989 17
rect 931 -51 989 -17
rect 931 -85 943 -51
rect 977 -85 989 -51
rect 931 -100 989 -85
<< pdiffc >>
rect -977 51 -943 85
rect -977 -17 -943 17
rect -977 -85 -943 -51
rect -849 51 -815 85
rect -849 -17 -815 17
rect -849 -85 -815 -51
rect -721 51 -687 85
rect -721 -17 -687 17
rect -721 -85 -687 -51
rect -593 51 -559 85
rect -593 -17 -559 17
rect -593 -85 -559 -51
rect -465 51 -431 85
rect -465 -17 -431 17
rect -465 -85 -431 -51
rect -337 51 -303 85
rect -337 -17 -303 17
rect -337 -85 -303 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -81 51 -47 85
rect -81 -17 -47 17
rect -81 -85 -47 -51
rect 47 51 81 85
rect 47 -17 81 17
rect 47 -85 81 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 303 51 337 85
rect 303 -17 337 17
rect 303 -85 337 -51
rect 431 51 465 85
rect 431 -17 465 17
rect 431 -85 465 -51
rect 559 51 593 85
rect 559 -17 593 17
rect 559 -85 593 -51
rect 687 51 721 85
rect 687 -17 721 17
rect 687 -85 721 -51
rect 815 51 849 85
rect 815 -17 849 17
rect 815 -85 849 -51
rect 943 51 977 85
rect 943 -17 977 17
rect 943 -85 977 -51
<< nsubdiff >>
rect -1091 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1091 283
rect -1091 187 -1057 249
rect -1091 119 -1057 153
rect 1057 187 1091 249
rect 1057 119 1091 153
rect -1091 51 -1057 85
rect -1091 -17 -1057 17
rect -1091 -85 -1057 -51
rect 1057 51 1091 85
rect 1057 -17 1091 17
rect 1057 -85 1091 -51
rect -1091 -153 -1057 -119
rect -1091 -249 -1057 -187
rect 1057 -153 1091 -119
rect 1057 -249 1091 -187
rect -1091 -283 -969 -249
rect -935 -283 -901 -249
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
rect 901 -283 935 -249
rect 969 -283 1091 -249
<< nsubdiffcont >>
rect -969 249 -935 283
rect -901 249 -867 283
rect -833 249 -799 283
rect -765 249 -731 283
rect -697 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 697 283
rect 731 249 765 283
rect 799 249 833 283
rect 867 249 901 283
rect 935 249 969 283
rect -1091 153 -1057 187
rect -1091 85 -1057 119
rect 1057 153 1091 187
rect -1091 17 -1057 51
rect -1091 -51 -1057 -17
rect -1091 -119 -1057 -85
rect 1057 85 1091 119
rect 1057 17 1091 51
rect 1057 -51 1091 -17
rect -1091 -187 -1057 -153
rect 1057 -119 1091 -85
rect 1057 -187 1091 -153
rect -969 -283 -935 -249
rect -901 -283 -867 -249
rect -833 -283 -799 -249
rect -765 -283 -731 -249
rect -697 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 697 -249
rect 731 -283 765 -249
rect 799 -283 833 -249
rect 867 -283 901 -249
rect 935 -283 969 -249
<< poly >>
rect -931 181 -861 197
rect -931 147 -913 181
rect -879 147 -861 181
rect -931 100 -861 147
rect -803 181 -733 197
rect -803 147 -785 181
rect -751 147 -733 181
rect -803 100 -733 147
rect -675 181 -605 197
rect -675 147 -657 181
rect -623 147 -605 181
rect -675 100 -605 147
rect -547 181 -477 197
rect -547 147 -529 181
rect -495 147 -477 181
rect -547 100 -477 147
rect -419 181 -349 197
rect -419 147 -401 181
rect -367 147 -349 181
rect -419 100 -349 147
rect -291 181 -221 197
rect -291 147 -273 181
rect -239 147 -221 181
rect -291 100 -221 147
rect -163 181 -93 197
rect -163 147 -145 181
rect -111 147 -93 181
rect -163 100 -93 147
rect -35 181 35 197
rect -35 147 -17 181
rect 17 147 35 181
rect -35 100 35 147
rect 93 181 163 197
rect 93 147 111 181
rect 145 147 163 181
rect 93 100 163 147
rect 221 181 291 197
rect 221 147 239 181
rect 273 147 291 181
rect 221 100 291 147
rect 349 181 419 197
rect 349 147 367 181
rect 401 147 419 181
rect 349 100 419 147
rect 477 181 547 197
rect 477 147 495 181
rect 529 147 547 181
rect 477 100 547 147
rect 605 181 675 197
rect 605 147 623 181
rect 657 147 675 181
rect 605 100 675 147
rect 733 181 803 197
rect 733 147 751 181
rect 785 147 803 181
rect 733 100 803 147
rect 861 181 931 197
rect 861 147 879 181
rect 913 147 931 181
rect 861 100 931 147
rect -931 -147 -861 -100
rect -931 -181 -913 -147
rect -879 -181 -861 -147
rect -931 -197 -861 -181
rect -803 -147 -733 -100
rect -803 -181 -785 -147
rect -751 -181 -733 -147
rect -803 -197 -733 -181
rect -675 -147 -605 -100
rect -675 -181 -657 -147
rect -623 -181 -605 -147
rect -675 -197 -605 -181
rect -547 -147 -477 -100
rect -547 -181 -529 -147
rect -495 -181 -477 -147
rect -547 -197 -477 -181
rect -419 -147 -349 -100
rect -419 -181 -401 -147
rect -367 -181 -349 -147
rect -419 -197 -349 -181
rect -291 -147 -221 -100
rect -291 -181 -273 -147
rect -239 -181 -221 -147
rect -291 -197 -221 -181
rect -163 -147 -93 -100
rect -163 -181 -145 -147
rect -111 -181 -93 -147
rect -163 -197 -93 -181
rect -35 -147 35 -100
rect -35 -181 -17 -147
rect 17 -181 35 -147
rect -35 -197 35 -181
rect 93 -147 163 -100
rect 93 -181 111 -147
rect 145 -181 163 -147
rect 93 -197 163 -181
rect 221 -147 291 -100
rect 221 -181 239 -147
rect 273 -181 291 -147
rect 221 -197 291 -181
rect 349 -147 419 -100
rect 349 -181 367 -147
rect 401 -181 419 -147
rect 349 -197 419 -181
rect 477 -147 547 -100
rect 477 -181 495 -147
rect 529 -181 547 -147
rect 477 -197 547 -181
rect 605 -147 675 -100
rect 605 -181 623 -147
rect 657 -181 675 -147
rect 605 -197 675 -181
rect 733 -147 803 -100
rect 733 -181 751 -147
rect 785 -181 803 -147
rect 733 -197 803 -181
rect 861 -147 931 -100
rect 861 -181 879 -147
rect 913 -181 931 -147
rect 861 -197 931 -181
<< polycont >>
rect -913 147 -879 181
rect -785 147 -751 181
rect -657 147 -623 181
rect -529 147 -495 181
rect -401 147 -367 181
rect -273 147 -239 181
rect -145 147 -111 181
rect -17 147 17 181
rect 111 147 145 181
rect 239 147 273 181
rect 367 147 401 181
rect 495 147 529 181
rect 623 147 657 181
rect 751 147 785 181
rect 879 147 913 181
rect -913 -181 -879 -147
rect -785 -181 -751 -147
rect -657 -181 -623 -147
rect -529 -181 -495 -147
rect -401 -181 -367 -147
rect -273 -181 -239 -147
rect -145 -181 -111 -147
rect -17 -181 17 -147
rect 111 -181 145 -147
rect 239 -181 273 -147
rect 367 -181 401 -147
rect 495 -181 529 -147
rect 623 -181 657 -147
rect 751 -181 785 -147
rect 879 -181 913 -147
<< locali >>
rect -1091 249 -969 283
rect -935 249 -901 283
rect -867 249 -833 283
rect -799 249 -765 283
rect -731 249 -697 283
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect 697 249 731 283
rect 765 249 799 283
rect 833 249 867 283
rect 901 249 935 283
rect 969 249 1091 283
rect -1091 187 -1057 249
rect 1057 187 1091 249
rect -1091 119 -1057 153
rect -931 147 -913 181
rect -879 147 -861 181
rect -803 147 -785 181
rect -751 147 -733 181
rect -675 147 -657 181
rect -623 147 -605 181
rect -547 147 -529 181
rect -495 147 -477 181
rect -419 147 -401 181
rect -367 147 -349 181
rect -291 147 -273 181
rect -239 147 -221 181
rect -163 147 -145 181
rect -111 147 -93 181
rect -35 147 -17 181
rect 17 147 35 181
rect 93 147 111 181
rect 145 147 163 181
rect 221 147 239 181
rect 273 147 291 181
rect 349 147 367 181
rect 401 147 419 181
rect 477 147 495 181
rect 529 147 547 181
rect 605 147 623 181
rect 657 147 675 181
rect 733 147 751 181
rect 785 147 803 181
rect 861 147 879 181
rect 913 147 931 181
rect 1057 119 1091 153
rect -1091 51 -1057 85
rect -1091 -17 -1057 17
rect -1091 -85 -1057 -51
rect -977 85 -943 104
rect -977 17 -943 19
rect -977 -19 -943 -17
rect -977 -104 -943 -85
rect -849 85 -815 104
rect -849 17 -815 19
rect -849 -19 -815 -17
rect -849 -104 -815 -85
rect -721 85 -687 104
rect -721 17 -687 19
rect -721 -19 -687 -17
rect -721 -104 -687 -85
rect -593 85 -559 104
rect -593 17 -559 19
rect -593 -19 -559 -17
rect -593 -104 -559 -85
rect -465 85 -431 104
rect -465 17 -431 19
rect -465 -19 -431 -17
rect -465 -104 -431 -85
rect -337 85 -303 104
rect -337 17 -303 19
rect -337 -19 -303 -17
rect -337 -104 -303 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -81 85 -47 104
rect -81 17 -47 19
rect -81 -19 -47 -17
rect -81 -104 -47 -85
rect 47 85 81 104
rect 47 17 81 19
rect 47 -19 81 -17
rect 47 -104 81 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 303 85 337 104
rect 303 17 337 19
rect 303 -19 337 -17
rect 303 -104 337 -85
rect 431 85 465 104
rect 431 17 465 19
rect 431 -19 465 -17
rect 431 -104 465 -85
rect 559 85 593 104
rect 559 17 593 19
rect 559 -19 593 -17
rect 559 -104 593 -85
rect 687 85 721 104
rect 687 17 721 19
rect 687 -19 721 -17
rect 687 -104 721 -85
rect 815 85 849 104
rect 815 17 849 19
rect 815 -19 849 -17
rect 815 -104 849 -85
rect 943 85 977 104
rect 943 17 977 19
rect 943 -19 977 -17
rect 943 -104 977 -85
rect 1057 51 1091 85
rect 1057 -17 1091 17
rect 1057 -85 1091 -51
rect -1091 -153 -1057 -119
rect -931 -181 -913 -147
rect -879 -181 -861 -147
rect -803 -181 -785 -147
rect -751 -181 -733 -147
rect -675 -181 -657 -147
rect -623 -181 -605 -147
rect -547 -181 -529 -147
rect -495 -181 -477 -147
rect -419 -181 -401 -147
rect -367 -181 -349 -147
rect -291 -181 -273 -147
rect -239 -181 -221 -147
rect -163 -181 -145 -147
rect -111 -181 -93 -147
rect -35 -181 -17 -147
rect 17 -181 35 -147
rect 93 -181 111 -147
rect 145 -181 163 -147
rect 221 -181 239 -147
rect 273 -181 291 -147
rect 349 -181 367 -147
rect 401 -181 419 -147
rect 477 -181 495 -147
rect 529 -181 547 -147
rect 605 -181 623 -147
rect 657 -181 675 -147
rect 733 -181 751 -147
rect 785 -181 803 -147
rect 861 -181 879 -147
rect 913 -181 931 -147
rect 1057 -153 1091 -119
rect -1091 -249 -1057 -187
rect 1057 -249 1091 -187
rect -1091 -283 -969 -249
rect -935 -283 -901 -249
rect -867 -283 -833 -249
rect -799 -283 -765 -249
rect -731 -283 -697 -249
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
rect 697 -283 731 -249
rect 765 -283 799 -249
rect 833 -283 867 -249
rect 901 -283 935 -249
rect 969 -283 1091 -249
<< viali >>
rect -913 147 -879 181
rect -785 147 -751 181
rect -657 147 -623 181
rect -529 147 -495 181
rect -401 147 -367 181
rect -273 147 -239 181
rect -145 147 -111 181
rect -17 147 17 181
rect 111 147 145 181
rect 239 147 273 181
rect 367 147 401 181
rect 495 147 529 181
rect 623 147 657 181
rect 751 147 785 181
rect 879 147 913 181
rect -977 51 -943 53
rect -977 19 -943 51
rect -977 -51 -943 -19
rect -977 -53 -943 -51
rect -849 51 -815 53
rect -849 19 -815 51
rect -849 -51 -815 -19
rect -849 -53 -815 -51
rect -721 51 -687 53
rect -721 19 -687 51
rect -721 -51 -687 -19
rect -721 -53 -687 -51
rect -593 51 -559 53
rect -593 19 -559 51
rect -593 -51 -559 -19
rect -593 -53 -559 -51
rect -465 51 -431 53
rect -465 19 -431 51
rect -465 -51 -431 -19
rect -465 -53 -431 -51
rect -337 51 -303 53
rect -337 19 -303 51
rect -337 -51 -303 -19
rect -337 -53 -303 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -81 51 -47 53
rect -81 19 -47 51
rect -81 -51 -47 -19
rect -81 -53 -47 -51
rect 47 51 81 53
rect 47 19 81 51
rect 47 -51 81 -19
rect 47 -53 81 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 303 51 337 53
rect 303 19 337 51
rect 303 -51 337 -19
rect 303 -53 337 -51
rect 431 51 465 53
rect 431 19 465 51
rect 431 -51 465 -19
rect 431 -53 465 -51
rect 559 51 593 53
rect 559 19 593 51
rect 559 -51 593 -19
rect 559 -53 593 -51
rect 687 51 721 53
rect 687 19 721 51
rect 687 -51 721 -19
rect 687 -53 721 -51
rect 815 51 849 53
rect 815 19 849 51
rect 815 -51 849 -19
rect 815 -53 849 -51
rect 943 51 977 53
rect 943 19 977 51
rect 943 -51 977 -19
rect 943 -53 977 -51
rect -913 -181 -879 -147
rect -785 -181 -751 -147
rect -657 -181 -623 -147
rect -529 -181 -495 -147
rect -401 -181 -367 -147
rect -273 -181 -239 -147
rect -145 -181 -111 -147
rect -17 -181 17 -147
rect 111 -181 145 -147
rect 239 -181 273 -147
rect 367 -181 401 -147
rect 495 -181 529 -147
rect 623 -181 657 -147
rect 751 -181 785 -147
rect 879 -181 913 -147
<< metal1 >>
rect -927 181 -865 187
rect -927 147 -913 181
rect -879 147 -865 181
rect -927 141 -865 147
rect -799 181 -737 187
rect -799 147 -785 181
rect -751 147 -737 181
rect -799 141 -737 147
rect -671 181 -609 187
rect -671 147 -657 181
rect -623 147 -609 181
rect -671 141 -609 147
rect -543 181 -481 187
rect -543 147 -529 181
rect -495 147 -481 181
rect -543 141 -481 147
rect -415 181 -353 187
rect -415 147 -401 181
rect -367 147 -353 181
rect -415 141 -353 147
rect -287 181 -225 187
rect -287 147 -273 181
rect -239 147 -225 181
rect -287 141 -225 147
rect -159 181 -97 187
rect -159 147 -145 181
rect -111 147 -97 181
rect -159 141 -97 147
rect -31 181 31 187
rect -31 147 -17 181
rect 17 147 31 181
rect -31 141 31 147
rect 97 181 159 187
rect 97 147 111 181
rect 145 147 159 181
rect 97 141 159 147
rect 225 181 287 187
rect 225 147 239 181
rect 273 147 287 181
rect 225 141 287 147
rect 353 181 415 187
rect 353 147 367 181
rect 401 147 415 181
rect 353 141 415 147
rect 481 181 543 187
rect 481 147 495 181
rect 529 147 543 181
rect 481 141 543 147
rect 609 181 671 187
rect 609 147 623 181
rect 657 147 671 181
rect 609 141 671 147
rect 737 181 799 187
rect 737 147 751 181
rect 785 147 799 181
rect 737 141 799 147
rect 865 181 927 187
rect 865 147 879 181
rect 913 147 927 181
rect 865 141 927 147
rect -983 53 -937 100
rect -983 19 -977 53
rect -943 19 -937 53
rect -983 -19 -937 19
rect -983 -53 -977 -19
rect -943 -53 -937 -19
rect -983 -100 -937 -53
rect -855 53 -809 100
rect -855 19 -849 53
rect -815 19 -809 53
rect -855 -19 -809 19
rect -855 -53 -849 -19
rect -815 -53 -809 -19
rect -855 -100 -809 -53
rect -727 53 -681 100
rect -727 19 -721 53
rect -687 19 -681 53
rect -727 -19 -681 19
rect -727 -53 -721 -19
rect -687 -53 -681 -19
rect -727 -100 -681 -53
rect -599 53 -553 100
rect -599 19 -593 53
rect -559 19 -553 53
rect -599 -19 -553 19
rect -599 -53 -593 -19
rect -559 -53 -553 -19
rect -599 -100 -553 -53
rect -471 53 -425 100
rect -471 19 -465 53
rect -431 19 -425 53
rect -471 -19 -425 19
rect -471 -53 -465 -19
rect -431 -53 -425 -19
rect -471 -100 -425 -53
rect -343 53 -297 100
rect -343 19 -337 53
rect -303 19 -297 53
rect -343 -19 -297 19
rect -343 -53 -337 -19
rect -303 -53 -297 -19
rect -343 -100 -297 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -87 53 -41 100
rect -87 19 -81 53
rect -47 19 -41 53
rect -87 -19 -41 19
rect -87 -53 -81 -19
rect -47 -53 -41 -19
rect -87 -100 -41 -53
rect 41 53 87 100
rect 41 19 47 53
rect 81 19 87 53
rect 41 -19 87 19
rect 41 -53 47 -19
rect 81 -53 87 -19
rect 41 -100 87 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 297 53 343 100
rect 297 19 303 53
rect 337 19 343 53
rect 297 -19 343 19
rect 297 -53 303 -19
rect 337 -53 343 -19
rect 297 -100 343 -53
rect 425 53 471 100
rect 425 19 431 53
rect 465 19 471 53
rect 425 -19 471 19
rect 425 -53 431 -19
rect 465 -53 471 -19
rect 425 -100 471 -53
rect 553 53 599 100
rect 553 19 559 53
rect 593 19 599 53
rect 553 -19 599 19
rect 553 -53 559 -19
rect 593 -53 599 -19
rect 553 -100 599 -53
rect 681 53 727 100
rect 681 19 687 53
rect 721 19 727 53
rect 681 -19 727 19
rect 681 -53 687 -19
rect 721 -53 727 -19
rect 681 -100 727 -53
rect 809 53 855 100
rect 809 19 815 53
rect 849 19 855 53
rect 809 -19 855 19
rect 809 -53 815 -19
rect 849 -53 855 -19
rect 809 -100 855 -53
rect 937 53 983 100
rect 937 19 943 53
rect 977 19 983 53
rect 937 -19 983 19
rect 937 -53 943 -19
rect 977 -53 983 -19
rect 937 -100 983 -53
rect -927 -147 -865 -141
rect -927 -181 -913 -147
rect -879 -181 -865 -147
rect -927 -187 -865 -181
rect -799 -147 -737 -141
rect -799 -181 -785 -147
rect -751 -181 -737 -147
rect -799 -187 -737 -181
rect -671 -147 -609 -141
rect -671 -181 -657 -147
rect -623 -181 -609 -147
rect -671 -187 -609 -181
rect -543 -147 -481 -141
rect -543 -181 -529 -147
rect -495 -181 -481 -147
rect -543 -187 -481 -181
rect -415 -147 -353 -141
rect -415 -181 -401 -147
rect -367 -181 -353 -147
rect -415 -187 -353 -181
rect -287 -147 -225 -141
rect -287 -181 -273 -147
rect -239 -181 -225 -147
rect -287 -187 -225 -181
rect -159 -147 -97 -141
rect -159 -181 -145 -147
rect -111 -181 -97 -147
rect -159 -187 -97 -181
rect -31 -147 31 -141
rect -31 -181 -17 -147
rect 17 -181 31 -147
rect -31 -187 31 -181
rect 97 -147 159 -141
rect 97 -181 111 -147
rect 145 -181 159 -147
rect 97 -187 159 -181
rect 225 -147 287 -141
rect 225 -181 239 -147
rect 273 -181 287 -147
rect 225 -187 287 -181
rect 353 -147 415 -141
rect 353 -181 367 -147
rect 401 -181 415 -147
rect 353 -187 415 -181
rect 481 -147 543 -141
rect 481 -181 495 -147
rect 529 -181 543 -147
rect 481 -187 543 -181
rect 609 -147 671 -141
rect 609 -181 623 -147
rect 657 -181 671 -147
rect 609 -187 671 -181
rect 737 -147 799 -141
rect 737 -181 751 -147
rect 785 -181 799 -147
rect 737 -187 799 -181
rect 865 -147 927 -141
rect 865 -181 879 -147
rect 913 -181 927 -147
rect 865 -187 927 -181
<< properties >>
string FIXED_BBOX -1074 -266 1074 266
<< end >>
