magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -812 -466 812 466
<< pmoslvt >>
rect -616 118 -416 318
rect -358 118 -158 318
rect -100 118 100 318
rect 158 118 358 318
rect 416 118 616 318
rect -616 -247 -416 -47
rect -358 -247 -158 -47
rect -100 -247 100 -47
rect 158 -247 358 -47
rect 416 -247 616 -47
<< pdiff >>
rect -674 303 -616 318
rect -674 269 -662 303
rect -628 269 -616 303
rect -674 235 -616 269
rect -674 201 -662 235
rect -628 201 -616 235
rect -674 167 -616 201
rect -674 133 -662 167
rect -628 133 -616 167
rect -674 118 -616 133
rect -416 303 -358 318
rect -416 269 -404 303
rect -370 269 -358 303
rect -416 235 -358 269
rect -416 201 -404 235
rect -370 201 -358 235
rect -416 167 -358 201
rect -416 133 -404 167
rect -370 133 -358 167
rect -416 118 -358 133
rect -158 303 -100 318
rect -158 269 -146 303
rect -112 269 -100 303
rect -158 235 -100 269
rect -158 201 -146 235
rect -112 201 -100 235
rect -158 167 -100 201
rect -158 133 -146 167
rect -112 133 -100 167
rect -158 118 -100 133
rect 100 303 158 318
rect 100 269 112 303
rect 146 269 158 303
rect 100 235 158 269
rect 100 201 112 235
rect 146 201 158 235
rect 100 167 158 201
rect 100 133 112 167
rect 146 133 158 167
rect 100 118 158 133
rect 358 303 416 318
rect 358 269 370 303
rect 404 269 416 303
rect 358 235 416 269
rect 358 201 370 235
rect 404 201 416 235
rect 358 167 416 201
rect 358 133 370 167
rect 404 133 416 167
rect 358 118 416 133
rect 616 303 674 318
rect 616 269 628 303
rect 662 269 674 303
rect 616 235 674 269
rect 616 201 628 235
rect 662 201 674 235
rect 616 167 674 201
rect 616 133 628 167
rect 662 133 674 167
rect 616 118 674 133
rect -674 -62 -616 -47
rect -674 -96 -662 -62
rect -628 -96 -616 -62
rect -674 -130 -616 -96
rect -674 -164 -662 -130
rect -628 -164 -616 -130
rect -674 -198 -616 -164
rect -674 -232 -662 -198
rect -628 -232 -616 -198
rect -674 -247 -616 -232
rect -416 -62 -358 -47
rect -416 -96 -404 -62
rect -370 -96 -358 -62
rect -416 -130 -358 -96
rect -416 -164 -404 -130
rect -370 -164 -358 -130
rect -416 -198 -358 -164
rect -416 -232 -404 -198
rect -370 -232 -358 -198
rect -416 -247 -358 -232
rect -158 -62 -100 -47
rect -158 -96 -146 -62
rect -112 -96 -100 -62
rect -158 -130 -100 -96
rect -158 -164 -146 -130
rect -112 -164 -100 -130
rect -158 -198 -100 -164
rect -158 -232 -146 -198
rect -112 -232 -100 -198
rect -158 -247 -100 -232
rect 100 -62 158 -47
rect 100 -96 112 -62
rect 146 -96 158 -62
rect 100 -130 158 -96
rect 100 -164 112 -130
rect 146 -164 158 -130
rect 100 -198 158 -164
rect 100 -232 112 -198
rect 146 -232 158 -198
rect 100 -247 158 -232
rect 358 -62 416 -47
rect 358 -96 370 -62
rect 404 -96 416 -62
rect 358 -130 416 -96
rect 358 -164 370 -130
rect 404 -164 416 -130
rect 358 -198 416 -164
rect 358 -232 370 -198
rect 404 -232 416 -198
rect 358 -247 416 -232
rect 616 -62 674 -47
rect 616 -96 628 -62
rect 662 -96 674 -62
rect 616 -130 674 -96
rect 616 -164 628 -130
rect 662 -164 674 -130
rect 616 -198 674 -164
rect 616 -232 628 -198
rect 662 -232 674 -198
rect 616 -247 674 -232
<< pdiffc >>
rect -662 269 -628 303
rect -662 201 -628 235
rect -662 133 -628 167
rect -404 269 -370 303
rect -404 201 -370 235
rect -404 133 -370 167
rect -146 269 -112 303
rect -146 201 -112 235
rect -146 133 -112 167
rect 112 269 146 303
rect 112 201 146 235
rect 112 133 146 167
rect 370 269 404 303
rect 370 201 404 235
rect 370 133 404 167
rect 628 269 662 303
rect 628 201 662 235
rect 628 133 662 167
rect -662 -96 -628 -62
rect -662 -164 -628 -130
rect -662 -232 -628 -198
rect -404 -96 -370 -62
rect -404 -164 -370 -130
rect -404 -232 -370 -198
rect -146 -96 -112 -62
rect -146 -164 -112 -130
rect -146 -232 -112 -198
rect 112 -96 146 -62
rect 112 -164 146 -130
rect 112 -232 146 -198
rect 370 -96 404 -62
rect 370 -164 404 -130
rect 370 -232 404 -198
rect 628 -96 662 -62
rect 628 -164 662 -130
rect 628 -232 662 -198
<< nsubdiff >>
rect -776 396 776 430
rect -776 -396 -742 396
rect 742 323 776 396
rect 742 255 776 289
rect 742 187 776 221
rect 742 119 776 153
rect 742 51 776 85
rect 742 -17 776 17
rect 742 -85 776 -51
rect 742 -153 776 -119
rect 742 -221 776 -187
rect 742 -289 776 -255
rect 742 -396 776 -323
rect -776 -430 776 -396
<< nsubdiffcont >>
rect 742 289 776 323
rect 742 221 776 255
rect 742 153 776 187
rect 742 85 776 119
rect 742 17 776 51
rect 742 -51 776 -17
rect 742 -119 776 -85
rect 742 -187 776 -153
rect 742 -255 776 -221
rect 742 -323 776 -289
<< poly >>
rect -616 318 -416 344
rect -358 318 -158 344
rect -100 318 100 344
rect 158 318 358 344
rect 416 318 616 344
rect -616 71 -416 118
rect -616 37 -567 71
rect -533 37 -499 71
rect -465 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -309 71
rect -275 37 -241 71
rect -207 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -51 71
rect -17 37 17 71
rect 51 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 207 71
rect 241 37 275 71
rect 309 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 465 71
rect 499 37 533 71
rect 567 37 616 71
rect 416 21 616 37
rect -616 -47 -416 -21
rect -358 -47 -158 -21
rect -100 -47 100 -21
rect 158 -47 358 -21
rect 416 -47 616 -21
rect -616 -294 -416 -247
rect -616 -328 -567 -294
rect -533 -328 -499 -294
rect -465 -328 -416 -294
rect -616 -344 -416 -328
rect -358 -294 -158 -247
rect -358 -328 -309 -294
rect -275 -328 -241 -294
rect -207 -328 -158 -294
rect -358 -344 -158 -328
rect -100 -294 100 -247
rect -100 -328 -51 -294
rect -17 -328 17 -294
rect 51 -328 100 -294
rect -100 -344 100 -328
rect 158 -294 358 -247
rect 158 -328 207 -294
rect 241 -328 275 -294
rect 309 -328 358 -294
rect 158 -344 358 -328
rect 416 -294 616 -247
rect 416 -328 465 -294
rect 499 -328 533 -294
rect 567 -328 616 -294
rect 416 -344 616 -328
<< polycont >>
rect -567 37 -533 71
rect -499 37 -465 71
rect -309 37 -275 71
rect -241 37 -207 71
rect -51 37 -17 71
rect 17 37 51 71
rect 207 37 241 71
rect 275 37 309 71
rect 465 37 499 71
rect 533 37 567 71
rect -567 -328 -533 -294
rect -499 -328 -465 -294
rect -309 -328 -275 -294
rect -241 -328 -207 -294
rect -51 -328 -17 -294
rect 17 -328 51 -294
rect 207 -328 241 -294
rect 275 -328 309 -294
rect 465 -328 499 -294
rect 533 -328 567 -294
<< locali >>
rect -776 396 776 430
rect -776 -396 -742 396
rect 742 323 776 396
rect -662 303 -628 322
rect -662 235 -628 237
rect -662 199 -628 201
rect -662 114 -628 133
rect -404 303 -370 322
rect -404 235 -370 237
rect -404 199 -370 201
rect -404 114 -370 133
rect -146 303 -112 322
rect -146 235 -112 237
rect -146 199 -112 201
rect -146 114 -112 133
rect 112 303 146 322
rect 112 235 146 237
rect 112 199 146 201
rect 112 114 146 133
rect 370 303 404 322
rect 370 235 404 237
rect 370 199 404 201
rect 370 114 404 133
rect 628 303 662 322
rect 628 235 662 237
rect 628 199 662 201
rect 628 114 662 133
rect 742 255 776 289
rect 742 187 776 221
rect 742 119 776 153
rect -616 37 -569 71
rect -533 37 -499 71
rect -463 37 -416 71
rect -358 37 -311 71
rect -275 37 -241 71
rect -205 37 -158 71
rect -100 37 -53 71
rect -17 37 17 71
rect 53 37 100 71
rect 158 37 205 71
rect 241 37 275 71
rect 311 37 358 71
rect 416 37 463 71
rect 499 37 533 71
rect 569 37 616 71
rect 742 51 776 85
rect 742 -17 776 17
rect -662 -62 -628 -43
rect -662 -130 -628 -128
rect -662 -166 -628 -164
rect -662 -251 -628 -232
rect -404 -62 -370 -43
rect -404 -130 -370 -128
rect -404 -166 -370 -164
rect -404 -251 -370 -232
rect -146 -62 -112 -43
rect -146 -130 -112 -128
rect -146 -166 -112 -164
rect -146 -251 -112 -232
rect 112 -62 146 -43
rect 112 -130 146 -128
rect 112 -166 146 -164
rect 112 -251 146 -232
rect 370 -62 404 -43
rect 370 -130 404 -128
rect 370 -166 404 -164
rect 370 -251 404 -232
rect 628 -62 662 -43
rect 628 -130 662 -128
rect 628 -166 662 -164
rect 628 -251 662 -232
rect 742 -85 776 -51
rect 742 -153 776 -119
rect 742 -221 776 -187
rect 742 -289 776 -255
rect -616 -328 -569 -294
rect -533 -328 -499 -294
rect -463 -328 -416 -294
rect -358 -328 -311 -294
rect -275 -328 -241 -294
rect -205 -328 -158 -294
rect -100 -328 -53 -294
rect -17 -328 17 -294
rect 53 -328 100 -294
rect 158 -328 205 -294
rect 241 -328 275 -294
rect 311 -328 358 -294
rect 416 -328 463 -294
rect 499 -328 533 -294
rect 569 -328 616 -294
rect 742 -396 776 -323
rect -776 -430 776 -396
<< viali >>
rect -662 269 -628 271
rect -662 237 -628 269
rect -662 167 -628 199
rect -662 165 -628 167
rect -404 269 -370 271
rect -404 237 -370 269
rect -404 167 -370 199
rect -404 165 -370 167
rect -146 269 -112 271
rect -146 237 -112 269
rect -146 167 -112 199
rect -146 165 -112 167
rect 112 269 146 271
rect 112 237 146 269
rect 112 167 146 199
rect 112 165 146 167
rect 370 269 404 271
rect 370 237 404 269
rect 370 167 404 199
rect 370 165 404 167
rect 628 269 662 271
rect 628 237 662 269
rect 628 167 662 199
rect 628 165 662 167
rect -569 37 -567 71
rect -567 37 -535 71
rect -497 37 -465 71
rect -465 37 -463 71
rect -311 37 -309 71
rect -309 37 -277 71
rect -239 37 -207 71
rect -207 37 -205 71
rect -53 37 -51 71
rect -51 37 -19 71
rect 19 37 51 71
rect 51 37 53 71
rect 205 37 207 71
rect 207 37 239 71
rect 277 37 309 71
rect 309 37 311 71
rect 463 37 465 71
rect 465 37 497 71
rect 535 37 567 71
rect 567 37 569 71
rect -662 -96 -628 -94
rect -662 -128 -628 -96
rect -662 -198 -628 -166
rect -662 -200 -628 -198
rect -404 -96 -370 -94
rect -404 -128 -370 -96
rect -404 -198 -370 -166
rect -404 -200 -370 -198
rect -146 -96 -112 -94
rect -146 -128 -112 -96
rect -146 -198 -112 -166
rect -146 -200 -112 -198
rect 112 -96 146 -94
rect 112 -128 146 -96
rect 112 -198 146 -166
rect 112 -200 146 -198
rect 370 -96 404 -94
rect 370 -128 404 -96
rect 370 -198 404 -166
rect 370 -200 404 -198
rect 628 -96 662 -94
rect 628 -128 662 -96
rect 628 -198 662 -166
rect 628 -200 662 -198
rect -569 -328 -567 -294
rect -567 -328 -535 -294
rect -497 -328 -465 -294
rect -465 -328 -463 -294
rect -311 -328 -309 -294
rect -309 -328 -277 -294
rect -239 -328 -207 -294
rect -207 -328 -205 -294
rect -53 -328 -51 -294
rect -51 -328 -19 -294
rect 19 -328 51 -294
rect 51 -328 53 -294
rect 205 -328 207 -294
rect 207 -328 239 -294
rect 277 -328 309 -294
rect 309 -328 311 -294
rect 463 -328 465 -294
rect 465 -328 497 -294
rect 535 -328 567 -294
rect 567 -328 569 -294
<< metal1 >>
rect -668 271 -622 318
rect -668 237 -662 271
rect -628 237 -622 271
rect -668 199 -622 237
rect -668 165 -662 199
rect -628 165 -622 199
rect -668 118 -622 165
rect -410 271 -364 318
rect -410 237 -404 271
rect -370 237 -364 271
rect -410 199 -364 237
rect -410 165 -404 199
rect -370 165 -364 199
rect -410 118 -364 165
rect -152 271 -106 318
rect -152 237 -146 271
rect -112 237 -106 271
rect -152 199 -106 237
rect -152 165 -146 199
rect -112 165 -106 199
rect -152 118 -106 165
rect 106 271 152 318
rect 106 237 112 271
rect 146 237 152 271
rect 106 199 152 237
rect 106 165 112 199
rect 146 165 152 199
rect 106 118 152 165
rect 364 271 410 318
rect 364 237 370 271
rect 404 237 410 271
rect 364 199 410 237
rect 364 165 370 199
rect 404 165 410 199
rect 364 118 410 165
rect 622 271 668 318
rect 622 237 628 271
rect 662 237 668 271
rect 622 199 668 237
rect 622 165 628 199
rect 662 165 668 199
rect 622 118 668 165
rect -612 71 -420 77
rect -612 37 -569 71
rect -535 37 -497 71
rect -463 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -311 71
rect -277 37 -239 71
rect -205 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -53 71
rect -19 37 19 71
rect 53 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 205 71
rect 239 37 277 71
rect 311 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 463 71
rect 497 37 535 71
rect 569 37 612 71
rect 420 31 612 37
rect -668 -94 -622 -47
rect -668 -128 -662 -94
rect -628 -128 -622 -94
rect -668 -166 -622 -128
rect -668 -200 -662 -166
rect -628 -200 -622 -166
rect -668 -247 -622 -200
rect -410 -94 -364 -47
rect -410 -128 -404 -94
rect -370 -128 -364 -94
rect -410 -166 -364 -128
rect -410 -200 -404 -166
rect -370 -200 -364 -166
rect -410 -247 -364 -200
rect -152 -94 -106 -47
rect -152 -128 -146 -94
rect -112 -128 -106 -94
rect -152 -166 -106 -128
rect -152 -200 -146 -166
rect -112 -200 -106 -166
rect -152 -247 -106 -200
rect 106 -94 152 -47
rect 106 -128 112 -94
rect 146 -128 152 -94
rect 106 -166 152 -128
rect 106 -200 112 -166
rect 146 -200 152 -166
rect 106 -247 152 -200
rect 364 -94 410 -47
rect 364 -128 370 -94
rect 404 -128 410 -94
rect 364 -166 410 -128
rect 364 -200 370 -166
rect 404 -200 410 -166
rect 364 -247 410 -200
rect 622 -94 668 -47
rect 622 -128 628 -94
rect 662 -128 668 -94
rect 622 -166 668 -128
rect 622 -200 628 -166
rect 662 -200 668 -166
rect 622 -247 668 -200
rect -612 -294 -420 -288
rect -612 -328 -569 -294
rect -535 -328 -497 -294
rect -463 -328 -420 -294
rect -612 -334 -420 -328
rect -354 -294 -162 -288
rect -354 -328 -311 -294
rect -277 -328 -239 -294
rect -205 -328 -162 -294
rect -354 -334 -162 -328
rect -96 -294 96 -288
rect -96 -328 -53 -294
rect -19 -328 19 -294
rect 53 -328 96 -294
rect -96 -334 96 -328
rect 162 -294 354 -288
rect 162 -328 205 -294
rect 239 -328 277 -294
rect 311 -328 354 -294
rect 162 -334 354 -328
rect 420 -294 612 -288
rect 420 -328 463 -294
rect 497 -328 535 -294
rect 569 -328 612 -294
rect 420 -334 612 -328
<< properties >>
string FIXED_BBOX -759 -413 759 413
<< end >>
