magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 3915 3945 4040 3980
rect 3265 3645 3380 3680
rect 4580 3650 4730 3685
rect 3260 3335 3385 3370
rect 3920 3335 4045 3370
rect 4580 3335 4705 3370
rect 3260 3185 3385 3220
rect 3890 3185 4070 3220
rect 4550 3185 4705 3220
rect 2435 2260 2470 2460
rect 3265 1035 3390 1070
rect 3920 1035 4045 1070
rect 4580 1035 4705 1070
<< metal1 >>
rect 3550 3881 3635 3900
rect 3550 3829 3566 3881
rect 3618 3829 3635 3881
rect 4325 3881 4410 3900
rect 3640 3868 3750 3874
rect 3738 3834 3750 3868
rect 3550 3810 3635 3829
rect 3640 3828 3750 3834
rect 3780 3831 3875 3845
rect 3665 3781 3750 3800
rect 3665 3778 3681 3781
rect 3550 3772 3681 3778
rect 3425 3731 3520 3745
rect 3550 3738 3562 3772
rect 3665 3738 3681 3772
rect 3550 3732 3681 3738
rect 3425 3679 3436 3731
rect 3488 3679 3520 3731
rect 3665 3729 3681 3732
rect 3733 3729 3750 3781
rect 3780 3779 3811 3831
rect 3863 3779 3875 3831
rect 3780 3765 3875 3779
rect 4085 3831 4180 3845
rect 4085 3779 4096 3831
rect 4148 3779 4180 3831
rect 4325 3829 4341 3881
rect 4393 3829 4410 3881
rect 4325 3810 4410 3829
rect 4085 3765 4180 3779
rect 4210 3781 4295 3800
rect 3665 3710 3750 3729
rect 4210 3729 4226 3781
rect 4278 3729 4295 3781
rect 4210 3710 4295 3729
rect 4440 3731 4535 3745
rect 3425 3665 3520 3679
rect 3550 3683 3635 3700
rect 3550 3631 3566 3683
rect 3618 3682 3635 3683
rect 4325 3683 4410 3700
rect 3618 3676 3750 3682
rect 3618 3642 3635 3676
rect 3738 3642 3750 3676
rect 3618 3636 3750 3642
rect 3780 3636 3875 3650
rect 3618 3631 3635 3636
rect 3550 3615 3635 3631
rect 3665 3588 3750 3605
rect 3665 3586 3681 3588
rect 3550 3580 3681 3586
rect 3425 3541 3520 3555
rect 2585 3521 3115 3530
rect 2585 3149 2600 3521
rect 3100 3149 3115 3521
rect 3425 3489 3436 3541
rect 3488 3489 3520 3541
rect 3550 3546 3562 3580
rect 3665 3546 3681 3580
rect 3550 3540 3681 3546
rect 3665 3536 3681 3540
rect 3733 3536 3750 3588
rect 3780 3584 3811 3636
rect 3863 3584 3875 3636
rect 3780 3570 3875 3584
rect 4085 3636 4180 3650
rect 4085 3584 4096 3636
rect 4148 3584 4180 3636
rect 4325 3631 4341 3683
rect 4393 3631 4410 3683
rect 4440 3679 4471 3731
rect 4523 3679 4535 3731
rect 4440 3665 4535 3679
rect 4325 3615 4410 3631
rect 4085 3570 4180 3584
rect 4210 3588 4295 3605
rect 3665 3520 3750 3536
rect 4210 3536 4226 3588
rect 4278 3536 4295 3588
rect 4210 3520 4295 3536
rect 4440 3541 4535 3555
rect 3425 3475 3520 3489
rect 3550 3491 3635 3510
rect 3550 3439 3566 3491
rect 3618 3490 3635 3491
rect 4325 3491 4410 3510
rect 3618 3484 3750 3490
rect 3618 3450 3635 3484
rect 3738 3450 3750 3484
rect 3618 3444 3750 3450
rect 3618 3439 3635 3444
rect 3550 3420 3635 3439
rect 4325 3439 4341 3491
rect 4393 3439 4410 3491
rect 4440 3489 4471 3541
rect 4523 3489 4535 3541
rect 4440 3475 4535 3489
rect 4845 3521 5375 3530
rect 4325 3420 4410 3439
rect 2585 3140 3115 3149
rect 4845 3149 4860 3521
rect 5360 3149 5375 3521
rect 4845 3140 5375 3149
rect 3665 3118 3750 3135
rect 3665 3110 3681 3118
rect 3550 3103 3681 3110
rect 3550 3070 3562 3103
rect 3665 3070 3681 3103
rect 3550 3066 3681 3070
rect 3733 3066 3750 3118
rect 4210 3118 4295 3135
rect 3550 3063 3750 3066
rect 3665 3050 3750 3063
rect 3780 3066 3875 3080
rect 3550 3018 3635 3035
rect 3425 2966 3520 2980
rect 3425 2914 3436 2966
rect 3488 2914 3520 2966
rect 3550 2966 3566 3018
rect 3618 3014 3635 3018
rect 3780 3014 3811 3066
rect 3863 3014 3875 3066
rect 3618 3007 3750 3014
rect 3618 2974 3635 3007
rect 3738 2974 3750 3007
rect 3780 3000 3875 3014
rect 4085 3066 4180 3080
rect 4085 3014 4096 3066
rect 4148 3014 4180 3066
rect 4210 3066 4226 3118
rect 4278 3110 4295 3118
rect 4278 3103 4410 3110
rect 4278 3070 4295 3103
rect 4398 3070 4410 3103
rect 4278 3066 4410 3070
rect 4210 3063 4410 3066
rect 4210 3050 4295 3063
rect 4325 3018 4410 3035
rect 4325 3014 4341 3018
rect 4085 3000 4180 3014
rect 4210 3007 4341 3014
rect 3618 2967 3750 2974
rect 4210 2974 4222 3007
rect 4325 2974 4341 3007
rect 4210 2967 4341 2974
rect 3618 2966 3635 2967
rect 3550 2950 3635 2966
rect 4325 2966 4341 2967
rect 4393 2966 4410 3018
rect 4325 2950 4410 2966
rect 4440 2966 4535 2980
rect 3665 2918 3750 2935
rect 3425 2900 3520 2914
rect 3550 2911 3681 2918
rect 3550 2878 3562 2911
rect 3665 2878 3681 2911
rect 3550 2871 3681 2878
rect 3665 2866 3681 2871
rect 3733 2866 3750 2918
rect 4210 2918 4295 2935
rect 3665 2850 3750 2866
rect 3780 2871 3875 2885
rect 3550 2823 3635 2840
rect 3425 2776 3520 2790
rect 3425 2724 3436 2776
rect 3488 2724 3520 2776
rect 3550 2771 3566 2823
rect 3618 2822 3635 2823
rect 3618 2815 3750 2822
rect 3618 2782 3635 2815
rect 3738 2782 3750 2815
rect 3780 2819 3811 2871
rect 3863 2819 3875 2871
rect 3780 2805 3875 2819
rect 4085 2871 4180 2885
rect 4085 2819 4096 2871
rect 4148 2819 4180 2871
rect 4210 2866 4226 2918
rect 4278 2911 4410 2918
rect 4278 2878 4295 2911
rect 4398 2878 4410 2911
rect 4440 2914 4471 2966
rect 4523 2914 4535 2966
rect 4440 2900 4535 2914
rect 4278 2871 4410 2878
rect 4278 2866 4295 2871
rect 4210 2850 4295 2866
rect 4325 2823 4410 2840
rect 4325 2822 4341 2823
rect 4085 2805 4180 2819
rect 4210 2815 4341 2822
rect 3618 2775 3750 2782
rect 4210 2782 4222 2815
rect 4325 2782 4341 2815
rect 4210 2775 4341 2782
rect 3618 2771 3635 2775
rect 3550 2755 3635 2771
rect 4325 2771 4341 2775
rect 4393 2771 4410 2823
rect 4325 2755 4410 2771
rect 4440 2776 4535 2790
rect 3665 2731 3750 2745
rect 3665 2726 3681 2731
rect 3425 2710 3520 2724
rect 3550 2718 3681 2726
rect 3550 2686 3562 2718
rect 3665 2686 3681 2718
rect 3550 2679 3681 2686
rect 3733 2679 3750 2731
rect 4210 2731 4295 2745
rect 3550 2678 3750 2679
rect 3665 2665 3750 2678
rect 3780 2681 3875 2695
rect 3550 2633 3635 2650
rect 3425 2586 3520 2600
rect 3425 2534 3436 2586
rect 3488 2534 3520 2586
rect 3550 2581 3566 2633
rect 3618 2630 3635 2633
rect 3618 2622 3750 2630
rect 3618 2590 3635 2622
rect 3738 2590 3750 2622
rect 3780 2629 3811 2681
rect 3863 2629 3875 2681
rect 3780 2615 3875 2629
rect 4085 2681 4180 2695
rect 4085 2629 4096 2681
rect 4148 2629 4180 2681
rect 4210 2679 4226 2731
rect 4278 2726 4295 2731
rect 4278 2718 4410 2726
rect 4278 2686 4295 2718
rect 4398 2686 4410 2718
rect 4440 2724 4471 2776
rect 4523 2724 4535 2776
rect 4440 2710 4535 2724
rect 4278 2679 4410 2686
rect 4210 2678 4410 2679
rect 4210 2665 4295 2678
rect 4325 2633 4410 2650
rect 4325 2630 4341 2633
rect 4085 2615 4180 2629
rect 4210 2622 4341 2630
rect 3618 2582 3750 2590
rect 4210 2590 4222 2622
rect 4325 2590 4341 2622
rect 4210 2582 4341 2590
rect 3618 2581 3635 2582
rect 3550 2565 3635 2581
rect 4325 2581 4341 2582
rect 4393 2581 4410 2633
rect 4325 2565 4410 2581
rect 4440 2586 4535 2600
rect 3665 2536 3750 2550
rect 3665 2534 3681 2536
rect 3425 2520 3520 2534
rect 3550 2526 3681 2534
rect 3550 2494 3562 2526
rect 3665 2494 3681 2526
rect 3550 2486 3681 2494
rect 3665 2484 3681 2486
rect 3733 2484 3750 2536
rect 4210 2536 4295 2550
rect 3665 2470 3750 2484
rect 3780 2486 3875 2500
rect 3550 2441 3635 2455
rect 3425 2396 3520 2410
rect 3425 2344 3436 2396
rect 3488 2344 3520 2396
rect 3550 2389 3566 2441
rect 3618 2438 3635 2441
rect 3618 2430 3750 2438
rect 3618 2398 3635 2430
rect 3738 2398 3750 2430
rect 3780 2434 3811 2486
rect 3863 2434 3875 2486
rect 3780 2420 3875 2434
rect 4085 2486 4180 2500
rect 4085 2434 4096 2486
rect 4148 2434 4180 2486
rect 4210 2484 4226 2536
rect 4278 2534 4295 2536
rect 4440 2534 4471 2586
rect 4523 2534 4535 2586
rect 4278 2526 4410 2534
rect 4278 2494 4295 2526
rect 4398 2494 4410 2526
rect 4440 2520 4535 2534
rect 4278 2486 4410 2494
rect 4278 2484 4295 2486
rect 4210 2470 4295 2484
rect 4325 2441 4410 2455
rect 4325 2438 4341 2441
rect 4085 2420 4180 2434
rect 4210 2430 4341 2438
rect 3618 2390 3750 2398
rect 4210 2398 4222 2430
rect 4325 2398 4341 2430
rect 4210 2390 4341 2398
rect 3618 2389 3635 2390
rect 3550 2375 3635 2389
rect 4325 2389 4341 2390
rect 4393 2389 4410 2441
rect 4325 2375 4410 2389
rect 4440 2396 4535 2410
rect 3665 2346 3750 2360
rect 3665 2344 3681 2346
rect 3425 2330 3520 2344
rect 3550 2336 3681 2344
rect 3550 2304 3562 2336
rect 3665 2304 3681 2336
rect 3550 2296 3681 2304
rect 3665 2294 3681 2296
rect 3733 2294 3750 2346
rect 4210 2346 4295 2360
rect 3665 2280 3750 2294
rect 3780 2296 3875 2310
rect 3550 2248 3635 2265
rect 3425 2201 3520 2215
rect 3425 2149 3436 2201
rect 3488 2149 3520 2201
rect 3550 2196 3566 2248
rect 3618 2240 3750 2248
rect 3618 2208 3635 2240
rect 3738 2208 3750 2240
rect 3780 2244 3811 2296
rect 3863 2244 3875 2296
rect 3780 2230 3875 2244
rect 4085 2296 4180 2310
rect 4085 2244 4096 2296
rect 4148 2244 4180 2296
rect 4210 2294 4226 2346
rect 4278 2344 4295 2346
rect 4440 2344 4471 2396
rect 4523 2344 4535 2396
rect 4278 2336 4410 2344
rect 4278 2304 4295 2336
rect 4398 2304 4410 2336
rect 4440 2330 4535 2344
rect 4278 2296 4410 2304
rect 4278 2294 4295 2296
rect 4210 2280 4295 2294
rect 4325 2248 4410 2265
rect 4085 2230 4180 2244
rect 4210 2240 4341 2248
rect 3618 2200 3750 2208
rect 4210 2208 4222 2240
rect 4325 2208 4341 2240
rect 4210 2200 4341 2208
rect 3618 2196 3635 2200
rect 3550 2180 3635 2196
rect 4325 2196 4341 2200
rect 4393 2196 4410 2248
rect 4325 2180 4410 2196
rect 4440 2201 4535 2215
rect 3665 2153 3750 2170
rect 3665 2152 3681 2153
rect 3425 2135 3520 2149
rect 3550 2144 3681 2152
rect 3550 2112 3562 2144
rect 3665 2112 3681 2144
rect 3550 2104 3681 2112
rect 3665 2101 3681 2104
rect 3733 2101 3750 2153
rect 4210 2153 4295 2170
rect 3665 2085 3750 2101
rect 3780 2106 3875 2120
rect 3550 2058 3635 2075
rect 3425 2011 3520 2025
rect 3425 1959 3436 2011
rect 3488 1959 3520 2011
rect 3550 2006 3566 2058
rect 3618 2056 3635 2058
rect 3618 2048 3750 2056
rect 3618 2016 3635 2048
rect 3738 2016 3750 2048
rect 3780 2054 3811 2106
rect 3863 2054 3875 2106
rect 3780 2040 3875 2054
rect 4085 2106 4180 2120
rect 4085 2054 4096 2106
rect 4148 2054 4180 2106
rect 4210 2101 4226 2153
rect 4278 2152 4295 2153
rect 4278 2144 4410 2152
rect 4278 2112 4295 2144
rect 4398 2112 4410 2144
rect 4440 2149 4471 2201
rect 4523 2149 4535 2201
rect 4440 2135 4535 2149
rect 4278 2104 4410 2112
rect 4278 2101 4295 2104
rect 4210 2085 4295 2101
rect 4325 2058 4410 2075
rect 4325 2056 4341 2058
rect 4085 2040 4180 2054
rect 4210 2048 4341 2056
rect 3618 2008 3750 2016
rect 4210 2016 4222 2048
rect 4325 2016 4341 2048
rect 4210 2008 4341 2016
rect 3618 2006 3635 2008
rect 3550 1990 3635 2006
rect 4325 2006 4341 2008
rect 4393 2006 4410 2058
rect 4325 1990 4410 2006
rect 4440 2011 4535 2025
rect 3665 1963 3750 1980
rect 3665 1959 3681 1963
rect 3425 1945 3520 1959
rect 3550 1952 3681 1959
rect 3550 1919 3562 1952
rect 3665 1919 3681 1952
rect 3550 1912 3681 1919
rect 3665 1911 3681 1912
rect 3733 1911 3750 1963
rect 4210 1963 4295 1980
rect 3665 1895 3750 1911
rect 3780 1911 3875 1925
rect 3550 1863 3635 1880
rect 3425 1816 3520 1830
rect 3425 1764 3436 1816
rect 3488 1764 3520 1816
rect 3550 1811 3566 1863
rect 3618 1856 3750 1863
rect 3618 1823 3635 1856
rect 3738 1823 3750 1856
rect 3780 1859 3811 1911
rect 3863 1859 3875 1911
rect 3780 1845 3875 1859
rect 4085 1911 4180 1925
rect 4085 1859 4096 1911
rect 4148 1859 4180 1911
rect 4210 1911 4226 1963
rect 4278 1959 4295 1963
rect 4440 1959 4471 2011
rect 4523 1959 4535 2011
rect 4278 1952 4410 1959
rect 4278 1919 4295 1952
rect 4398 1919 4410 1952
rect 4440 1945 4535 1959
rect 4278 1912 4410 1919
rect 4278 1911 4295 1912
rect 4210 1895 4295 1911
rect 4325 1863 4410 1880
rect 4085 1845 4180 1859
rect 4210 1856 4341 1863
rect 3618 1816 3750 1823
rect 4210 1823 4222 1856
rect 4325 1823 4341 1856
rect 4210 1816 4341 1823
rect 3618 1811 3635 1816
rect 3550 1795 3635 1811
rect 4325 1811 4341 1816
rect 4393 1811 4410 1863
rect 4325 1795 4410 1811
rect 4440 1816 4535 1830
rect 3665 1768 3750 1785
rect 3665 1767 3681 1768
rect 3425 1750 3520 1764
rect 3550 1760 3681 1767
rect 3550 1727 3562 1760
rect 3665 1727 3681 1760
rect 3550 1720 3681 1727
rect 3665 1716 3681 1720
rect 3733 1716 3750 1768
rect 4210 1768 4295 1785
rect 3665 1700 3750 1716
rect 3780 1721 3875 1735
rect 3550 1673 3635 1690
rect 3425 1626 3520 1640
rect 2565 1568 3135 1600
rect 2565 1196 2600 1568
rect 3100 1196 3135 1568
rect 3425 1574 3436 1626
rect 3488 1574 3520 1626
rect 3550 1621 3566 1673
rect 3618 1671 3635 1673
rect 3618 1664 3750 1671
rect 3618 1631 3635 1664
rect 3738 1631 3750 1664
rect 3780 1669 3811 1721
rect 3863 1669 3875 1721
rect 3780 1655 3875 1669
rect 4085 1721 4180 1735
rect 4085 1669 4096 1721
rect 4148 1669 4180 1721
rect 4210 1716 4226 1768
rect 4278 1767 4295 1768
rect 4278 1760 4410 1767
rect 4278 1727 4295 1760
rect 4398 1727 4410 1760
rect 4440 1764 4471 1816
rect 4523 1764 4535 1816
rect 4440 1750 4535 1764
rect 4278 1720 4410 1727
rect 4278 1716 4295 1720
rect 4210 1700 4295 1716
rect 4325 1673 4410 1690
rect 4325 1671 4341 1673
rect 4085 1655 4180 1669
rect 4210 1664 4341 1671
rect 3618 1624 3750 1631
rect 4210 1631 4222 1664
rect 4325 1631 4341 1664
rect 4210 1624 4341 1631
rect 3618 1621 3635 1624
rect 3550 1605 3635 1621
rect 4325 1621 4341 1624
rect 4393 1621 4410 1673
rect 4325 1605 4410 1621
rect 4440 1626 4535 1640
rect 3665 1578 3750 1595
rect 3665 1574 3681 1578
rect 3425 1560 3520 1574
rect 3550 1568 3681 1574
rect 3550 1534 3562 1568
rect 3665 1534 3681 1568
rect 3550 1528 3681 1534
rect 3665 1526 3681 1528
rect 3733 1526 3750 1578
rect 4210 1578 4295 1595
rect 3665 1510 3750 1526
rect 3780 1526 3875 1540
rect 3550 1478 3635 1500
rect 3425 1431 3520 1445
rect 3425 1379 3436 1431
rect 3488 1379 3520 1431
rect 3550 1426 3566 1478
rect 3618 1472 3750 1478
rect 3618 1438 3635 1472
rect 3738 1438 3750 1472
rect 3780 1474 3811 1526
rect 3863 1474 3875 1526
rect 3780 1460 3875 1474
rect 4085 1526 4180 1540
rect 4085 1474 4096 1526
rect 4148 1474 4180 1526
rect 4210 1526 4226 1578
rect 4278 1574 4295 1578
rect 4440 1574 4471 1626
rect 4523 1574 4535 1626
rect 4278 1568 4410 1574
rect 4278 1534 4295 1568
rect 4398 1534 4410 1568
rect 4440 1560 4535 1574
rect 4825 1568 5395 1600
rect 4278 1528 4410 1534
rect 4278 1526 4295 1528
rect 4210 1510 4295 1526
rect 4325 1478 4410 1500
rect 4085 1460 4180 1474
rect 4210 1472 4341 1478
rect 3618 1432 3750 1438
rect 4210 1438 4222 1472
rect 4325 1438 4341 1472
rect 4210 1432 4341 1438
rect 3618 1426 3635 1432
rect 3550 1410 3635 1426
rect 4325 1426 4341 1432
rect 4393 1426 4410 1478
rect 4325 1410 4410 1426
rect 4440 1431 4535 1445
rect 3665 1383 3750 1400
rect 3665 1382 3681 1383
rect 3425 1365 3520 1379
rect 3550 1376 3681 1382
rect 3550 1342 3562 1376
rect 3665 1342 3681 1376
rect 3550 1336 3681 1342
rect 3665 1331 3681 1336
rect 3733 1331 3750 1383
rect 4210 1383 4295 1400
rect 3665 1315 3750 1331
rect 3780 1336 3875 1350
rect 3550 1288 3635 1305
rect 2565 1165 3135 1196
rect 3425 1241 3520 1255
rect 3425 1189 3436 1241
rect 3488 1189 3520 1241
rect 3550 1236 3566 1288
rect 3618 1286 3635 1288
rect 3618 1280 3750 1286
rect 3618 1246 3635 1280
rect 3738 1246 3750 1280
rect 3780 1284 3811 1336
rect 3863 1284 3875 1336
rect 3780 1270 3875 1284
rect 4085 1336 4180 1350
rect 4085 1284 4096 1336
rect 4148 1284 4180 1336
rect 4210 1331 4226 1383
rect 4278 1382 4295 1383
rect 4278 1376 4410 1382
rect 4278 1342 4295 1376
rect 4398 1342 4410 1376
rect 4440 1379 4471 1431
rect 4523 1379 4535 1431
rect 4440 1365 4535 1379
rect 4278 1336 4410 1342
rect 4278 1331 4295 1336
rect 4210 1315 4295 1331
rect 4325 1288 4410 1305
rect 4325 1286 4341 1288
rect 4085 1270 4180 1284
rect 4210 1280 4341 1286
rect 3618 1240 3750 1246
rect 4210 1246 4222 1280
rect 4325 1246 4341 1280
rect 4210 1240 4341 1246
rect 3618 1236 3635 1240
rect 3550 1220 3635 1236
rect 4325 1236 4341 1240
rect 4393 1236 4410 1288
rect 4325 1220 4410 1236
rect 4440 1241 4535 1255
rect 3665 1191 3750 1210
rect 3665 1190 3681 1191
rect 3425 1175 3520 1189
rect 3550 1184 3681 1190
rect 3550 1150 3562 1184
rect 3665 1150 3681 1184
rect 3550 1144 3681 1150
rect 3665 1139 3681 1144
rect 3733 1139 3750 1191
rect 3665 1120 3750 1139
rect 4210 1191 4295 1210
rect 4210 1139 4226 1191
rect 4278 1190 4295 1191
rect 4278 1184 4410 1190
rect 4278 1150 4295 1184
rect 4398 1150 4410 1184
rect 4440 1189 4471 1241
rect 4523 1189 4535 1241
rect 4440 1175 4535 1189
rect 4825 1196 4860 1568
rect 5360 1196 5395 1568
rect 4825 1165 5395 1196
rect 4278 1144 4410 1150
rect 4278 1139 4295 1144
rect 4210 1120 4295 1139
<< via1 >>
rect 3566 3829 3618 3881
rect 3436 3679 3488 3731
rect 3681 3729 3733 3781
rect 3811 3779 3863 3831
rect 4096 3779 4148 3831
rect 4341 3829 4393 3881
rect 4226 3729 4278 3781
rect 3566 3631 3618 3683
rect 2600 3149 3100 3521
rect 3436 3489 3488 3541
rect 3681 3536 3733 3588
rect 3811 3584 3863 3636
rect 4096 3584 4148 3636
rect 4341 3631 4393 3683
rect 4471 3679 4523 3731
rect 4226 3536 4278 3588
rect 3566 3439 3618 3491
rect 4341 3439 4393 3491
rect 4471 3489 4523 3541
rect 4860 3149 5360 3521
rect 3681 3066 3733 3118
rect 3436 2914 3488 2966
rect 3566 2966 3618 3018
rect 3811 3014 3863 3066
rect 4096 3014 4148 3066
rect 4226 3066 4278 3118
rect 4341 2966 4393 3018
rect 3681 2866 3733 2918
rect 3436 2724 3488 2776
rect 3566 2771 3618 2823
rect 3811 2819 3863 2871
rect 4096 2819 4148 2871
rect 4226 2866 4278 2918
rect 4471 2914 4523 2966
rect 4341 2771 4393 2823
rect 3681 2679 3733 2731
rect 3436 2534 3488 2586
rect 3566 2581 3618 2633
rect 3811 2629 3863 2681
rect 4096 2629 4148 2681
rect 4226 2679 4278 2731
rect 4471 2724 4523 2776
rect 4341 2581 4393 2633
rect 3681 2484 3733 2536
rect 3436 2344 3488 2396
rect 3566 2389 3618 2441
rect 3811 2434 3863 2486
rect 4096 2434 4148 2486
rect 4226 2484 4278 2536
rect 4471 2534 4523 2586
rect 4341 2389 4393 2441
rect 3681 2294 3733 2346
rect 3436 2149 3488 2201
rect 3566 2196 3618 2248
rect 3811 2244 3863 2296
rect 4096 2244 4148 2296
rect 4226 2294 4278 2346
rect 4471 2344 4523 2396
rect 4341 2196 4393 2248
rect 3681 2101 3733 2153
rect 3436 1959 3488 2011
rect 3566 2006 3618 2058
rect 3811 2054 3863 2106
rect 4096 2054 4148 2106
rect 4226 2101 4278 2153
rect 4471 2149 4523 2201
rect 4341 2006 4393 2058
rect 3681 1911 3733 1963
rect 3436 1764 3488 1816
rect 3566 1811 3618 1863
rect 3811 1859 3863 1911
rect 4096 1859 4148 1911
rect 4226 1911 4278 1963
rect 4471 1959 4523 2011
rect 4341 1811 4393 1863
rect 3681 1716 3733 1768
rect 2600 1196 3100 1568
rect 3436 1574 3488 1626
rect 3566 1621 3618 1673
rect 3811 1669 3863 1721
rect 4096 1669 4148 1721
rect 4226 1716 4278 1768
rect 4471 1764 4523 1816
rect 4341 1621 4393 1673
rect 3681 1526 3733 1578
rect 3436 1379 3488 1431
rect 3566 1426 3618 1478
rect 3811 1474 3863 1526
rect 4096 1474 4148 1526
rect 4226 1526 4278 1578
rect 4471 1574 4523 1626
rect 4341 1426 4393 1478
rect 3681 1331 3733 1383
rect 3436 1189 3488 1241
rect 3566 1236 3618 1288
rect 3811 1284 3863 1336
rect 4096 1284 4148 1336
rect 4226 1331 4278 1383
rect 4471 1379 4523 1431
rect 4341 1236 4393 1288
rect 3681 1139 3733 1191
rect 4226 1139 4278 1191
rect 4471 1189 4523 1241
rect 4860 1196 5360 1568
<< metal2 >>
rect 3425 3945 3875 4020
rect 3425 3731 3500 3945
rect 3530 3883 3635 3900
rect 3530 3827 3547 3883
rect 3603 3881 3635 3883
rect 3618 3829 3635 3881
rect 3603 3827 3635 3829
rect 3530 3810 3635 3827
rect 3800 3831 3875 3945
rect 3425 3679 3436 3731
rect 3488 3679 3500 3731
rect 3665 3783 3770 3800
rect 3665 3781 3697 3783
rect 3665 3729 3681 3781
rect 3665 3727 3697 3729
rect 3753 3727 3770 3783
rect 3665 3710 3770 3727
rect 3800 3779 3811 3831
rect 3863 3779 3875 3831
rect 2565 3523 3135 3550
rect 2565 3521 2622 3523
rect 3078 3521 3135 3523
rect 2565 3149 2600 3521
rect 3100 3149 3135 3521
rect 3425 3541 3500 3679
rect 3530 3685 3635 3700
rect 3530 3629 3547 3685
rect 3603 3683 3635 3685
rect 3618 3631 3635 3683
rect 3603 3629 3635 3631
rect 3530 3615 3635 3629
rect 3800 3636 3875 3779
rect 3425 3489 3436 3541
rect 3488 3489 3500 3541
rect 3665 3590 3770 3605
rect 3665 3588 3697 3590
rect 3665 3536 3681 3588
rect 3665 3534 3697 3536
rect 3753 3534 3770 3590
rect 3800 3584 3811 3636
rect 3863 3584 3875 3636
rect 3800 3570 3875 3584
rect 4085 3945 4535 4020
rect 4085 3831 4160 3945
rect 4085 3779 4096 3831
rect 4148 3779 4160 3831
rect 4325 3883 4430 3900
rect 4325 3881 4357 3883
rect 4325 3829 4341 3881
rect 4325 3827 4357 3829
rect 4413 3827 4430 3883
rect 4325 3810 4430 3827
rect 4085 3636 4160 3779
rect 4190 3783 4295 3800
rect 4190 3727 4207 3783
rect 4263 3781 4295 3783
rect 4278 3729 4295 3781
rect 4263 3727 4295 3729
rect 4190 3710 4295 3727
rect 4460 3731 4535 3945
rect 4085 3584 4096 3636
rect 4148 3584 4160 3636
rect 4325 3685 4430 3700
rect 4325 3683 4357 3685
rect 4325 3631 4341 3683
rect 4325 3629 4357 3631
rect 4413 3629 4430 3685
rect 4325 3615 4430 3629
rect 4460 3679 4471 3731
rect 4523 3679 4535 3731
rect 4085 3570 4160 3584
rect 4190 3590 4295 3605
rect 3665 3520 3770 3534
rect 4190 3534 4207 3590
rect 4263 3588 4295 3590
rect 4278 3536 4295 3588
rect 4263 3534 4295 3536
rect 4190 3520 4295 3534
rect 4460 3541 4535 3679
rect 3425 3475 3500 3489
rect 3530 3493 3635 3510
rect 3530 3437 3547 3493
rect 3603 3491 3635 3493
rect 3618 3439 3635 3491
rect 3603 3437 3635 3439
rect 3530 3420 3635 3437
rect 4325 3493 4430 3510
rect 4325 3491 4357 3493
rect 4325 3439 4341 3491
rect 4325 3437 4357 3439
rect 4413 3437 4430 3493
rect 4460 3489 4471 3541
rect 4523 3489 4535 3541
rect 4460 3475 4535 3489
rect 4825 3523 5395 3550
rect 4825 3521 4882 3523
rect 5338 3521 5395 3523
rect 4325 3420 4430 3437
rect 2565 3147 2622 3149
rect 3078 3147 3135 3149
rect 2565 3120 3135 3147
rect 4825 3149 4860 3521
rect 5360 3149 5395 3521
rect 4825 3147 4882 3149
rect 5338 3147 5395 3149
rect 3665 3120 3770 3135
rect 3665 3118 3697 3120
rect 3665 3066 3681 3118
rect 3665 3064 3697 3066
rect 3753 3064 3770 3120
rect 4190 3120 4295 3135
rect 4825 3120 5395 3147
rect 3665 3050 3770 3064
rect 3800 3066 3875 3080
rect 3535 3020 3635 3035
rect 3425 2966 3500 2980
rect 3425 2914 3436 2966
rect 3488 2914 3500 2966
rect 3535 2964 3547 3020
rect 3603 3018 3635 3020
rect 3618 2966 3635 3018
rect 3603 2964 3635 2966
rect 3535 2950 3635 2964
rect 3800 3014 3811 3066
rect 3863 3014 3875 3066
rect 3425 2776 3500 2914
rect 3665 2920 3770 2935
rect 3665 2918 3697 2920
rect 3665 2866 3681 2918
rect 3665 2864 3697 2866
rect 3753 2864 3770 2920
rect 3665 2850 3770 2864
rect 3800 2871 3875 3014
rect 3425 2724 3436 2776
rect 3488 2724 3500 2776
rect 3535 2825 3635 2840
rect 3535 2769 3547 2825
rect 3603 2823 3635 2825
rect 3618 2771 3635 2823
rect 3603 2769 3635 2771
rect 3535 2755 3635 2769
rect 3800 2819 3811 2871
rect 3863 2819 3875 2871
rect 3425 2586 3500 2724
rect 3665 2733 3770 2750
rect 3665 2731 3697 2733
rect 3665 2679 3681 2731
rect 3665 2677 3697 2679
rect 3753 2677 3770 2733
rect 3665 2665 3770 2677
rect 3800 2681 3875 2819
rect 3425 2534 3436 2586
rect 3488 2534 3500 2586
rect 3535 2635 3635 2650
rect 3535 2579 3547 2635
rect 3603 2633 3635 2635
rect 3618 2581 3635 2633
rect 3603 2579 3635 2581
rect 3535 2565 3635 2579
rect 3800 2629 3811 2681
rect 3863 2629 3875 2681
rect 3425 2396 3500 2534
rect 3665 2538 3770 2550
rect 3665 2536 3697 2538
rect 3665 2484 3681 2536
rect 3665 2482 3697 2484
rect 3753 2482 3770 2538
rect 3665 2470 3770 2482
rect 3800 2486 3875 2629
rect 3425 2344 3436 2396
rect 3488 2344 3500 2396
rect 3535 2443 3635 2455
rect 3535 2387 3547 2443
rect 3603 2441 3635 2443
rect 3618 2389 3635 2441
rect 3603 2387 3635 2389
rect 3535 2375 3635 2387
rect 3800 2434 3811 2486
rect 3863 2434 3875 2486
rect 3425 2201 3500 2344
rect 3665 2348 3770 2365
rect 3665 2346 3697 2348
rect 3665 2294 3681 2346
rect 3665 2292 3697 2294
rect 3753 2292 3770 2348
rect 3665 2280 3770 2292
rect 3800 2296 3875 2434
rect 3425 2149 3436 2201
rect 3488 2149 3500 2201
rect 3535 2250 3635 2265
rect 3535 2194 3547 2250
rect 3603 2248 3635 2250
rect 3618 2196 3635 2248
rect 3603 2194 3635 2196
rect 3535 2180 3635 2194
rect 3800 2244 3811 2296
rect 3863 2244 3875 2296
rect 3425 2011 3500 2149
rect 3665 2155 3770 2170
rect 3665 2153 3697 2155
rect 3665 2101 3681 2153
rect 3665 2099 3697 2101
rect 3753 2099 3770 2155
rect 3665 2085 3770 2099
rect 3800 2106 3875 2244
rect 3425 1959 3436 2011
rect 3488 1959 3500 2011
rect 3535 2060 3635 2075
rect 3535 2004 3547 2060
rect 3603 2058 3635 2060
rect 3618 2006 3635 2058
rect 3603 2004 3635 2006
rect 3535 1990 3635 2004
rect 3800 2054 3811 2106
rect 3863 2054 3875 2106
rect 3425 1816 3500 1959
rect 3665 1965 3770 1980
rect 3665 1963 3697 1965
rect 3665 1911 3681 1963
rect 3665 1909 3697 1911
rect 3753 1909 3770 1965
rect 3665 1895 3770 1909
rect 3800 1911 3875 2054
rect 3425 1764 3436 1816
rect 3488 1764 3500 1816
rect 3535 1865 3635 1880
rect 3535 1809 3547 1865
rect 3603 1863 3635 1865
rect 3618 1811 3635 1863
rect 3603 1809 3635 1811
rect 3535 1795 3635 1809
rect 3800 1859 3811 1911
rect 3863 1859 3875 1911
rect 3425 1626 3500 1764
rect 3665 1770 3770 1785
rect 3665 1768 3697 1770
rect 3665 1716 3681 1768
rect 3665 1714 3697 1716
rect 3753 1714 3770 1770
rect 3665 1700 3770 1714
rect 3800 1721 3875 1859
rect 2565 1568 3135 1600
rect 2565 1196 2600 1568
rect 3100 1196 3135 1568
rect 2565 590 3135 1196
rect 2565 374 2622 590
rect 3078 374 3135 590
rect 2565 335 3135 374
rect 3425 1574 3436 1626
rect 3488 1574 3500 1626
rect 3535 1675 3635 1690
rect 3535 1619 3547 1675
rect 3603 1673 3635 1675
rect 3618 1621 3635 1673
rect 3603 1619 3635 1621
rect 3535 1605 3635 1619
rect 3800 1669 3811 1721
rect 3863 1669 3875 1721
rect 3425 1431 3500 1574
rect 3665 1580 3770 1595
rect 3665 1578 3697 1580
rect 3665 1526 3681 1578
rect 3665 1524 3697 1526
rect 3753 1524 3770 1580
rect 3665 1510 3770 1524
rect 3800 1526 3875 1669
rect 3425 1379 3436 1431
rect 3488 1379 3500 1431
rect 3535 1480 3635 1495
rect 3535 1424 3547 1480
rect 3603 1478 3635 1480
rect 3618 1426 3635 1478
rect 3603 1424 3635 1426
rect 3535 1410 3635 1424
rect 3800 1474 3811 1526
rect 3863 1474 3875 1526
rect 3425 1241 3500 1379
rect 3665 1385 3770 1400
rect 3665 1383 3697 1385
rect 3665 1331 3681 1383
rect 3665 1329 3697 1331
rect 3753 1329 3770 1385
rect 3665 1315 3770 1329
rect 3800 1336 3875 1474
rect 3425 1189 3436 1241
rect 3488 1189 3500 1241
rect 3530 1290 3635 1305
rect 3530 1234 3547 1290
rect 3603 1288 3635 1290
rect 3618 1236 3635 1288
rect 3603 1234 3635 1236
rect 3530 1220 3635 1234
rect 3800 1284 3811 1336
rect 3863 1284 3875 1336
rect 3425 305 3500 1189
rect 3665 1193 3770 1210
rect 3665 1191 3697 1193
rect 3665 1139 3681 1191
rect 3665 1137 3697 1139
rect 3753 1137 3770 1193
rect 3665 1120 3770 1137
rect 3800 305 3875 1284
rect 4085 3066 4160 3080
rect 4085 3014 4096 3066
rect 4148 3014 4160 3066
rect 4190 3064 4207 3120
rect 4263 3118 4295 3120
rect 4278 3066 4295 3118
rect 4263 3064 4295 3066
rect 4190 3050 4295 3064
rect 4085 2871 4160 3014
rect 4325 3020 4425 3035
rect 4325 3018 4357 3020
rect 4325 2966 4341 3018
rect 4325 2964 4357 2966
rect 4413 2964 4425 3020
rect 4325 2950 4425 2964
rect 4460 2966 4535 2980
rect 4085 2819 4096 2871
rect 4148 2819 4160 2871
rect 4190 2920 4295 2935
rect 4190 2864 4207 2920
rect 4263 2918 4295 2920
rect 4278 2866 4295 2918
rect 4263 2864 4295 2866
rect 4190 2850 4295 2864
rect 4460 2914 4471 2966
rect 4523 2914 4535 2966
rect 4085 2681 4160 2819
rect 4325 2825 4425 2840
rect 4325 2823 4357 2825
rect 4325 2771 4341 2823
rect 4325 2769 4357 2771
rect 4413 2769 4425 2825
rect 4325 2755 4425 2769
rect 4460 2776 4535 2914
rect 4085 2629 4096 2681
rect 4148 2629 4160 2681
rect 4190 2733 4295 2750
rect 4190 2677 4207 2733
rect 4263 2731 4295 2733
rect 4278 2679 4295 2731
rect 4263 2677 4295 2679
rect 4190 2665 4295 2677
rect 4460 2724 4471 2776
rect 4523 2724 4535 2776
rect 4085 2486 4160 2629
rect 4325 2635 4425 2650
rect 4325 2633 4357 2635
rect 4325 2581 4341 2633
rect 4325 2579 4357 2581
rect 4413 2579 4425 2635
rect 4325 2565 4425 2579
rect 4460 2586 4535 2724
rect 4085 2434 4096 2486
rect 4148 2434 4160 2486
rect 4190 2538 4295 2550
rect 4190 2482 4207 2538
rect 4263 2536 4295 2538
rect 4278 2484 4295 2536
rect 4263 2482 4295 2484
rect 4190 2470 4295 2482
rect 4460 2534 4471 2586
rect 4523 2534 4535 2586
rect 4085 2296 4160 2434
rect 4325 2443 4425 2455
rect 4325 2441 4357 2443
rect 4325 2389 4341 2441
rect 4325 2387 4357 2389
rect 4413 2387 4425 2443
rect 4325 2375 4425 2387
rect 4460 2396 4535 2534
rect 4085 2244 4096 2296
rect 4148 2244 4160 2296
rect 4190 2348 4295 2365
rect 4190 2292 4207 2348
rect 4263 2346 4295 2348
rect 4278 2294 4295 2346
rect 4263 2292 4295 2294
rect 4190 2280 4295 2292
rect 4460 2344 4471 2396
rect 4523 2344 4535 2396
rect 4085 2106 4160 2244
rect 4325 2250 4425 2265
rect 4325 2248 4357 2250
rect 4325 2196 4341 2248
rect 4325 2194 4357 2196
rect 4413 2194 4425 2250
rect 4325 2180 4425 2194
rect 4460 2201 4535 2344
rect 4085 2054 4096 2106
rect 4148 2054 4160 2106
rect 4190 2155 4295 2170
rect 4190 2099 4207 2155
rect 4263 2153 4295 2155
rect 4278 2101 4295 2153
rect 4263 2099 4295 2101
rect 4190 2085 4295 2099
rect 4460 2149 4471 2201
rect 4523 2149 4535 2201
rect 4085 1911 4160 2054
rect 4325 2060 4425 2075
rect 4325 2058 4357 2060
rect 4325 2006 4341 2058
rect 4325 2004 4357 2006
rect 4413 2004 4425 2060
rect 4325 1990 4425 2004
rect 4460 2011 4535 2149
rect 4085 1859 4096 1911
rect 4148 1859 4160 1911
rect 4190 1965 4295 1980
rect 4190 1909 4207 1965
rect 4263 1963 4295 1965
rect 4278 1911 4295 1963
rect 4263 1909 4295 1911
rect 4190 1895 4295 1909
rect 4460 1959 4471 2011
rect 4523 1959 4535 2011
rect 4085 1721 4160 1859
rect 4325 1865 4425 1880
rect 4325 1863 4357 1865
rect 4325 1811 4341 1863
rect 4325 1809 4357 1811
rect 4413 1809 4425 1865
rect 4325 1795 4425 1809
rect 4460 1816 4535 1959
rect 4085 1669 4096 1721
rect 4148 1669 4160 1721
rect 4190 1770 4295 1785
rect 4190 1714 4207 1770
rect 4263 1768 4295 1770
rect 4278 1716 4295 1768
rect 4263 1714 4295 1716
rect 4190 1700 4295 1714
rect 4460 1764 4471 1816
rect 4523 1764 4535 1816
rect 4085 1526 4160 1669
rect 4325 1675 4425 1690
rect 4325 1673 4357 1675
rect 4325 1621 4341 1673
rect 4325 1619 4357 1621
rect 4413 1619 4425 1675
rect 4325 1605 4425 1619
rect 4460 1626 4535 1764
rect 4085 1474 4096 1526
rect 4148 1474 4160 1526
rect 4190 1580 4295 1595
rect 4190 1524 4207 1580
rect 4263 1578 4295 1580
rect 4278 1526 4295 1578
rect 4263 1524 4295 1526
rect 4190 1510 4295 1524
rect 4460 1574 4471 1626
rect 4523 1574 4535 1626
rect 4085 1336 4160 1474
rect 4325 1480 4425 1495
rect 4325 1478 4357 1480
rect 4325 1426 4341 1478
rect 4325 1424 4357 1426
rect 4413 1424 4425 1480
rect 4325 1410 4425 1424
rect 4460 1431 4535 1574
rect 4085 1284 4096 1336
rect 4148 1284 4160 1336
rect 4190 1385 4295 1400
rect 4190 1329 4207 1385
rect 4263 1383 4295 1385
rect 4278 1331 4295 1383
rect 4263 1329 4295 1331
rect 4190 1315 4295 1329
rect 4460 1379 4471 1431
rect 4523 1379 4535 1431
rect 4085 305 4160 1284
rect 4325 1290 4430 1305
rect 4325 1288 4357 1290
rect 4325 1236 4341 1288
rect 4325 1234 4357 1236
rect 4413 1234 4430 1290
rect 4325 1220 4430 1234
rect 4460 1241 4535 1379
rect 4190 1193 4295 1210
rect 4190 1137 4207 1193
rect 4263 1191 4295 1193
rect 4278 1139 4295 1191
rect 4263 1137 4295 1139
rect 4190 1120 4295 1137
rect 4460 1189 4471 1241
rect 4523 1189 4535 1241
rect 4460 305 4535 1189
rect 4825 1568 5395 1600
rect 4825 1196 4860 1568
rect 5360 1196 5395 1568
rect 4825 593 5395 1196
rect 4825 377 4882 593
rect 5338 377 5395 593
rect 4825 335 5395 377
rect 2400 230 4535 305
<< via2 >>
rect 3547 3881 3603 3883
rect 3547 3829 3566 3881
rect 3566 3829 3603 3881
rect 3547 3827 3603 3829
rect 3697 3781 3753 3783
rect 3697 3729 3733 3781
rect 3733 3729 3753 3781
rect 3697 3727 3753 3729
rect 2622 3521 3078 3523
rect 2622 3149 3078 3521
rect 3547 3683 3603 3685
rect 3547 3631 3566 3683
rect 3566 3631 3603 3683
rect 3547 3629 3603 3631
rect 3697 3588 3753 3590
rect 3697 3536 3733 3588
rect 3733 3536 3753 3588
rect 3697 3534 3753 3536
rect 4357 3881 4413 3883
rect 4357 3829 4393 3881
rect 4393 3829 4413 3881
rect 4357 3827 4413 3829
rect 4207 3781 4263 3783
rect 4207 3729 4226 3781
rect 4226 3729 4263 3781
rect 4207 3727 4263 3729
rect 4357 3683 4413 3685
rect 4357 3631 4393 3683
rect 4393 3631 4413 3683
rect 4357 3629 4413 3631
rect 4207 3588 4263 3590
rect 4207 3536 4226 3588
rect 4226 3536 4263 3588
rect 4207 3534 4263 3536
rect 3547 3491 3603 3493
rect 3547 3439 3566 3491
rect 3566 3439 3603 3491
rect 3547 3437 3603 3439
rect 4357 3491 4413 3493
rect 4357 3439 4393 3491
rect 4393 3439 4413 3491
rect 4357 3437 4413 3439
rect 4882 3521 5338 3523
rect 2622 3147 3078 3149
rect 4882 3149 5338 3521
rect 4882 3147 5338 3149
rect 3697 3118 3753 3120
rect 3697 3066 3733 3118
rect 3733 3066 3753 3118
rect 3697 3064 3753 3066
rect 3547 3018 3603 3020
rect 3547 2966 3566 3018
rect 3566 2966 3603 3018
rect 3547 2964 3603 2966
rect 3697 2918 3753 2920
rect 3697 2866 3733 2918
rect 3733 2866 3753 2918
rect 3697 2864 3753 2866
rect 3547 2823 3603 2825
rect 3547 2771 3566 2823
rect 3566 2771 3603 2823
rect 3547 2769 3603 2771
rect 3697 2731 3753 2733
rect 3697 2679 3733 2731
rect 3733 2679 3753 2731
rect 3697 2677 3753 2679
rect 3547 2633 3603 2635
rect 3547 2581 3566 2633
rect 3566 2581 3603 2633
rect 3547 2579 3603 2581
rect 3697 2536 3753 2538
rect 3697 2484 3733 2536
rect 3733 2484 3753 2536
rect 3697 2482 3753 2484
rect 3547 2441 3603 2443
rect 3547 2389 3566 2441
rect 3566 2389 3603 2441
rect 3547 2387 3603 2389
rect 3697 2346 3753 2348
rect 3697 2294 3733 2346
rect 3733 2294 3753 2346
rect 3697 2292 3753 2294
rect 3547 2248 3603 2250
rect 3547 2196 3566 2248
rect 3566 2196 3603 2248
rect 3547 2194 3603 2196
rect 3697 2153 3753 2155
rect 3697 2101 3733 2153
rect 3733 2101 3753 2153
rect 3697 2099 3753 2101
rect 3547 2058 3603 2060
rect 3547 2006 3566 2058
rect 3566 2006 3603 2058
rect 3547 2004 3603 2006
rect 3697 1963 3753 1965
rect 3697 1911 3733 1963
rect 3733 1911 3753 1963
rect 3697 1909 3753 1911
rect 3547 1863 3603 1865
rect 3547 1811 3566 1863
rect 3566 1811 3603 1863
rect 3547 1809 3603 1811
rect 3697 1768 3753 1770
rect 3697 1716 3733 1768
rect 3733 1716 3753 1768
rect 3697 1714 3753 1716
rect 2622 374 3078 590
rect 3547 1673 3603 1675
rect 3547 1621 3566 1673
rect 3566 1621 3603 1673
rect 3547 1619 3603 1621
rect 3697 1578 3753 1580
rect 3697 1526 3733 1578
rect 3733 1526 3753 1578
rect 3697 1524 3753 1526
rect 3547 1478 3603 1480
rect 3547 1426 3566 1478
rect 3566 1426 3603 1478
rect 3547 1424 3603 1426
rect 3697 1383 3753 1385
rect 3697 1331 3733 1383
rect 3733 1331 3753 1383
rect 3697 1329 3753 1331
rect 3547 1288 3603 1290
rect 3547 1236 3566 1288
rect 3566 1236 3603 1288
rect 3547 1234 3603 1236
rect 3697 1191 3753 1193
rect 3697 1139 3733 1191
rect 3733 1139 3753 1191
rect 3697 1137 3753 1139
rect 4207 3118 4263 3120
rect 4207 3066 4226 3118
rect 4226 3066 4263 3118
rect 4207 3064 4263 3066
rect 4357 3018 4413 3020
rect 4357 2966 4393 3018
rect 4393 2966 4413 3018
rect 4357 2964 4413 2966
rect 4207 2918 4263 2920
rect 4207 2866 4226 2918
rect 4226 2866 4263 2918
rect 4207 2864 4263 2866
rect 4357 2823 4413 2825
rect 4357 2771 4393 2823
rect 4393 2771 4413 2823
rect 4357 2769 4413 2771
rect 4207 2731 4263 2733
rect 4207 2679 4226 2731
rect 4226 2679 4263 2731
rect 4207 2677 4263 2679
rect 4357 2633 4413 2635
rect 4357 2581 4393 2633
rect 4393 2581 4413 2633
rect 4357 2579 4413 2581
rect 4207 2536 4263 2538
rect 4207 2484 4226 2536
rect 4226 2484 4263 2536
rect 4207 2482 4263 2484
rect 4357 2441 4413 2443
rect 4357 2389 4393 2441
rect 4393 2389 4413 2441
rect 4357 2387 4413 2389
rect 4207 2346 4263 2348
rect 4207 2294 4226 2346
rect 4226 2294 4263 2346
rect 4207 2292 4263 2294
rect 4357 2248 4413 2250
rect 4357 2196 4393 2248
rect 4393 2196 4413 2248
rect 4357 2194 4413 2196
rect 4207 2153 4263 2155
rect 4207 2101 4226 2153
rect 4226 2101 4263 2153
rect 4207 2099 4263 2101
rect 4357 2058 4413 2060
rect 4357 2006 4393 2058
rect 4393 2006 4413 2058
rect 4357 2004 4413 2006
rect 4207 1963 4263 1965
rect 4207 1911 4226 1963
rect 4226 1911 4263 1963
rect 4207 1909 4263 1911
rect 4357 1863 4413 1865
rect 4357 1811 4393 1863
rect 4393 1811 4413 1863
rect 4357 1809 4413 1811
rect 4207 1768 4263 1770
rect 4207 1716 4226 1768
rect 4226 1716 4263 1768
rect 4207 1714 4263 1716
rect 4357 1673 4413 1675
rect 4357 1621 4393 1673
rect 4393 1621 4413 1673
rect 4357 1619 4413 1621
rect 4207 1578 4263 1580
rect 4207 1526 4226 1578
rect 4226 1526 4263 1578
rect 4207 1524 4263 1526
rect 4357 1478 4413 1480
rect 4357 1426 4393 1478
rect 4393 1426 4413 1478
rect 4357 1424 4413 1426
rect 4207 1383 4263 1385
rect 4207 1331 4226 1383
rect 4226 1331 4263 1383
rect 4207 1329 4263 1331
rect 4357 1288 4413 1290
rect 4357 1236 4393 1288
rect 4393 1236 4413 1288
rect 4357 1234 4413 1236
rect 4207 1191 4263 1193
rect 4207 1139 4226 1191
rect 4226 1139 4263 1191
rect 4207 1137 4263 1139
rect 4882 377 5338 593
<< metal3 >>
rect 3320 3883 3620 3900
rect 3320 3827 3547 3883
rect 3603 3827 3620 3883
rect 4340 3883 4640 3900
rect 3320 3685 3620 3827
rect 3320 3629 3547 3685
rect 3603 3629 3620 3685
rect 3320 3600 3620 3629
rect 2566 3523 3620 3600
rect 2566 3147 2622 3523
rect 3078 3493 3620 3523
rect 3078 3437 3547 3493
rect 3603 3437 3620 3493
rect 3078 3300 3620 3437
rect 3680 3783 4280 3845
rect 3680 3727 3697 3783
rect 3753 3727 4207 3783
rect 4263 3727 4280 3783
rect 3680 3590 4280 3727
rect 3680 3534 3697 3590
rect 3753 3534 4207 3590
rect 4263 3534 4280 3590
rect 3078 3147 3135 3300
rect 2566 3120 3135 3147
rect 3680 3155 4280 3534
rect 4340 3827 4357 3883
rect 4413 3827 4640 3883
rect 4340 3685 4640 3827
rect 4340 3629 4357 3685
rect 4413 3629 4640 3685
rect 4340 3600 4640 3629
rect 4340 3550 5395 3600
rect 4340 3523 5396 3550
rect 4340 3493 4882 3523
rect 4340 3437 4357 3493
rect 4413 3437 4882 3493
rect 4340 3300 4882 3437
rect 3320 3020 3620 3140
rect 3320 2964 3547 3020
rect 3603 2964 3620 3020
rect 3320 2825 3620 2964
rect 3320 2769 3547 2825
rect 3603 2769 3620 2825
rect 3320 2635 3620 2769
rect 3320 2579 3547 2635
rect 3603 2579 3620 2635
rect 3320 2443 3620 2579
rect 3320 2387 3547 2443
rect 3603 2387 3620 2443
rect 3320 2250 3620 2387
rect 3320 2194 3547 2250
rect 3603 2194 3620 2250
rect 3320 2060 3620 2194
rect 3320 2004 3547 2060
rect 3603 2004 3620 2060
rect 3320 1865 3620 2004
rect 3320 1809 3547 1865
rect 3603 1809 3620 1865
rect 3320 1675 3620 1809
rect 3320 1619 3547 1675
rect 3603 1619 3620 1675
rect 3320 1480 3620 1619
rect 3320 1424 3547 1480
rect 3603 1424 3620 1480
rect 3320 1290 3620 1424
rect 3320 1234 3547 1290
rect 3603 1234 3620 1290
rect 3320 1045 3620 1234
rect 3680 3120 3800 3155
rect 3680 3064 3697 3120
rect 3753 3080 3800 3120
rect 3875 3120 4280 3155
rect 4825 3147 4882 3300
rect 5338 3147 5396 3523
rect 3875 3080 4207 3120
rect 3753 3064 4207 3080
rect 4263 3064 4280 3120
rect 3680 2920 4280 3064
rect 3680 2864 3697 2920
rect 3753 2864 4207 2920
rect 4263 2864 4280 2920
rect 3680 2733 4280 2864
rect 3680 2677 3697 2733
rect 3753 2677 4207 2733
rect 4263 2677 4280 2733
rect 3680 2538 4280 2677
rect 3680 2482 3697 2538
rect 3753 2482 4207 2538
rect 4263 2482 4280 2538
rect 3680 2348 4280 2482
rect 3680 2292 3697 2348
rect 3753 2292 4207 2348
rect 4263 2292 4280 2348
rect 3680 2155 4280 2292
rect 3680 2099 3697 2155
rect 3753 2099 4207 2155
rect 4263 2099 4280 2155
rect 3680 1965 4280 2099
rect 3680 1909 3697 1965
rect 3753 1909 4207 1965
rect 4263 1909 4280 1965
rect 3680 1770 4280 1909
rect 3680 1714 3697 1770
rect 3753 1714 4207 1770
rect 4263 1714 4280 1770
rect 3680 1580 4280 1714
rect 3680 1524 3697 1580
rect 3753 1524 4207 1580
rect 4263 1524 4280 1580
rect 3680 1385 4280 1524
rect 3680 1329 3697 1385
rect 3753 1329 4207 1385
rect 4263 1329 4280 1385
rect 3680 1193 4280 1329
rect 3680 1137 3697 1193
rect 3753 1137 4207 1193
rect 4263 1137 4280 1193
rect 3680 1105 4280 1137
rect 4340 3020 4640 3140
rect 4825 3120 5396 3147
rect 4340 2964 4357 3020
rect 4413 2964 4640 3020
rect 4340 2825 4640 2964
rect 4340 2769 4357 2825
rect 4413 2769 4640 2825
rect 4340 2635 4640 2769
rect 4340 2579 4357 2635
rect 4413 2579 4640 2635
rect 4340 2443 4640 2579
rect 4340 2387 4357 2443
rect 4413 2387 4640 2443
rect 4340 2250 4640 2387
rect 4340 2194 4357 2250
rect 4413 2194 4640 2250
rect 4340 2060 4640 2194
rect 4340 2004 4357 2060
rect 4413 2004 4640 2060
rect 4340 1865 4640 2004
rect 4340 1809 4357 1865
rect 4413 1809 4640 1865
rect 4340 1675 4640 1809
rect 4340 1619 4357 1675
rect 4413 1619 4640 1675
rect 4340 1480 4640 1619
rect 4340 1424 4357 1480
rect 4413 1424 4640 1480
rect 4340 1290 4640 1424
rect 4340 1234 4357 1290
rect 4413 1234 4640 1290
rect 4340 1045 4640 1234
rect 2400 745 4640 1045
rect 2400 695 2700 745
rect 2400 593 5395 635
rect 2400 590 4882 593
rect 2400 374 2622 590
rect 3078 377 4882 590
rect 5338 377 5395 593
rect 3078 374 5395 377
rect 2400 335 5395 374
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM1
timestamp 1663011646
transform 0 -1 3650 -1 0 2127
box -1117 -300 1117 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM2
timestamp 1663011646
transform 0 -1 3650 -1 0 3659
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM3
timestamp 1663011646
transform 0 1 4310 -1 0 3659
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM4
timestamp 1663011646
transform 0 1 4310 -1 0 2127
box -1117 -300 1117 300
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR16
timestamp 1663011646
transform 1 0 2851 0 1 2358
box -441 -1348 441 1348
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR17
timestamp 1663011646
transform 1 0 5111 0 1 2358
box -441 -1348 441 1348
<< labels >>
flabel metal2 s 3425 3945 3875 4020 1 FreeMono 2 0 0 0 INA
port 1 nsew
flabel metal2 s 4085 3945 4535 4020 1 FreeMono 2 0 0 0 INB
port 2 nsew
flabel metal3 s 2400 335 2585 635 1 FreeMono 2 0 0 0 VDD
port 3 nsew
flabel metal2 s 2400 230 4535 305 1 FreeMono 2 0 0 0 BIAS
port 4 nsew
rlabel metal2 s 2457 267 2457 267 4 BIAS
port 4 nsew
rlabel metal2 s 3467 267 3467 267 4 BIAS
port 4 nsew
rlabel metal3 s 2492 485 2492 485 4 VDD
port 3 nsew
rlabel metal3 s 2400 695 2700 1045 4 GND
port 5 nsew
rlabel metal2 s 3650 3982 3650 3982 4 INA
port 1 nsew
rlabel metal2 s 4310 3982 4310 3982 4 INB
port 2 nsew
rlabel locali s 2435 2260 2470 2460 4 SUB
port 6 nsew
rlabel metal3 s 2566 3552 3136 3598 4 OUTA
port 7 nsew
rlabel metal3 s 4340 3530 5395 3600 4 OUTB
port 8 nsew
<< end >>
