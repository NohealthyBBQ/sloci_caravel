magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal1 >>
rect 14920 682865 15420 682910
rect 14920 682045 14989 682865
rect 15361 682045 15420 682865
rect 14920 668280 15420 682045
rect 14920 668180 23410 668280
rect 14920 668100 23840 668180
rect 14920 668060 23410 668100
rect 55960 662576 56100 662620
rect 55960 662524 56004 662576
rect 56056 662524 56100 662576
rect 55960 662480 56100 662524
rect 56200 661656 56340 661700
rect 56200 661604 56244 661656
rect 56296 661604 56340 661656
rect 56200 661560 56340 661604
rect 56480 661056 56620 661100
rect 56480 661004 56524 661056
rect 56576 661004 56620 661056
rect 56480 660960 56620 661004
rect 56720 660536 56860 660580
rect 56720 660484 56764 660536
rect 56816 660484 56860 660536
rect 56720 660440 56860 660484
rect 56980 660176 57120 660220
rect 56980 660124 57024 660176
rect 57076 660124 57120 660176
rect 56980 660080 57120 660124
<< via1 >>
rect 14989 682045 15361 682865
rect 56004 662524 56056 662576
rect 56244 661604 56296 661656
rect 56524 661004 56576 661056
rect 56764 660484 56816 660536
rect 57024 660124 57076 660176
<< metal2 >>
rect 14920 682865 15420 682910
rect 14920 682843 14989 682865
rect 15361 682843 15420 682865
rect 14920 682067 14987 682843
rect 15363 682067 15420 682843
rect 14920 682045 14989 682067
rect 15361 682045 15420 682067
rect 14920 681990 15420 682045
rect 23190 671593 25400 671620
rect 23190 671457 23222 671593
rect 23358 671457 25400 671593
rect 23190 671420 25400 671457
rect 55960 662576 56100 662620
rect 55960 662524 56004 662576
rect 56056 662524 56100 662576
rect 55960 335218 56100 662524
rect 56200 661656 56340 661700
rect 56200 661604 56244 661656
rect 56296 661604 56340 661656
rect 56200 378458 56340 661604
rect 56480 661056 56620 661100
rect 56480 661004 56524 661056
rect 56576 661004 56620 661056
rect 56480 421658 56620 661004
rect 56720 660536 56860 660580
rect 56720 660484 56764 660536
rect 56816 660484 56860 660536
rect 56720 466078 56860 660484
rect 56980 660176 57120 660220
rect 56980 660124 57024 660176
rect 57076 660124 57120 660176
rect 56980 508118 57120 660124
rect 238000 590968 246800 592200
rect 238000 582032 239032 590968
rect 245968 582032 246800 590968
rect 238000 580200 246800 582032
rect 246300 579400 246700 580200
rect 56980 508062 57022 508118
rect 57078 508062 57120 508118
rect 56980 508038 57120 508062
rect 56980 507982 57022 508038
rect 57078 507982 57120 508038
rect 56980 507960 57120 507982
rect 56720 466022 56762 466078
rect 56818 466022 56860 466078
rect 56720 465998 56860 466022
rect 56720 465942 56762 465998
rect 56818 465942 56860 465998
rect 56720 465920 56860 465942
rect 56480 421602 56522 421658
rect 56578 421602 56620 421658
rect 56480 421578 56620 421602
rect 56480 421522 56522 421578
rect 56578 421522 56620 421578
rect 56480 421500 56620 421522
rect 56200 378402 56242 378458
rect 56298 378402 56340 378458
rect 56200 378378 56340 378402
rect 56200 378322 56242 378378
rect 56298 378322 56340 378378
rect 56200 378300 56340 378322
rect 55960 335162 56002 335218
rect 56058 335162 56100 335218
rect 55960 335138 56100 335162
rect 55960 335082 56002 335138
rect 56058 335082 56100 335138
rect 55960 335060 56100 335082
<< via2 >>
rect 14987 682067 14989 682843
rect 14989 682067 15361 682843
rect 15361 682067 15363 682843
rect 23222 671457 23358 671593
rect 239032 582032 245968 590968
rect 57022 508062 57078 508118
rect 57022 507982 57078 508038
rect 56762 466022 56818 466078
rect 56762 465942 56818 465998
rect 56522 421602 56578 421658
rect 56522 421522 56578 421578
rect 56242 378402 56298 378458
rect 56242 378322 56298 378378
rect 56002 335162 56058 335218
rect 56002 335082 56058 335138
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 703200 125194 704800
rect 17070 689360 19380 702300
rect 68470 689480 70760 702300
rect 42500 689437 70760 689480
rect 17070 689330 26050 689360
rect 17070 688210 41870 689330
rect 42500 688413 42598 689437
rect 43142 688413 70760 689437
rect 42500 688360 70760 688413
rect 120000 701000 125200 703200
rect 165594 702300 170594 704800
rect 173394 703000 175594 704800
rect 173394 702300 175600 703000
rect 175894 702300 180894 704800
rect 510594 703000 515394 704800
rect 520594 703000 525394 704800
rect 173400 701772 175600 702300
rect 17070 688200 26050 688210
rect -800 682910 1700 685242
rect -800 682843 15420 682910
rect -800 682067 14987 682843
rect 15363 682067 15420 682843
rect -800 681990 15420 682067
rect -800 680242 1700 681990
rect 40710 680350 41870 688210
rect 40720 679110 41870 680350
rect 40720 677237 41720 677320
rect 40720 676133 40773 677237
rect 41637 676133 41720 677237
rect 40720 676080 41720 676133
rect 23190 671593 23390 671620
rect 23190 671457 23222 671593
rect 23358 671457 23390 671593
rect 23190 669072 23390 671457
rect 23190 668688 23218 669072
rect 23362 668688 23390 669072
rect 23190 668640 23390 668688
rect -800 648600 1660 648642
rect -800 646992 80246 648600
rect -800 643842 73008 646992
rect 246 638642 73008 643842
rect -800 635008 73008 638642
rect 78992 635008 80246 646992
rect -800 633842 80246 635008
rect 246 633838 80246 633842
rect 120000 606000 124000 701000
rect 173400 699628 173628 701772
rect 175372 699628 175600 701772
rect 173400 699200 175600 699628
rect 510000 701992 526000 703000
rect 510000 694008 511008 701992
rect 524992 694008 526000 701992
rect 510000 693000 526000 694008
rect 570200 644584 583800 644600
rect 570200 642992 584800 644584
rect 570200 631008 572008 642992
rect 579992 639784 584800 642992
rect 579992 634584 583800 639784
rect 579992 631008 584800 634584
rect 570200 629800 584800 631008
rect 582340 629784 584800 629800
rect 21990 605992 24010 606000
rect 21990 604008 22008 605992
rect 23992 604008 24010 605992
rect 21990 604000 24010 604008
rect 22000 596000 24000 604000
rect 120000 602000 288000 606000
rect 22000 594000 285400 596000
rect 238990 591000 246010 591005
rect 164000 590968 246010 591000
rect 164000 589972 239032 590968
rect 164000 583028 165028 589972
rect 181972 583028 239032 589972
rect 164000 582032 239032 583028
rect 245968 582032 246010 590968
rect 164000 582000 246010 582032
rect 154000 581400 158000 582000
rect 238990 581995 246010 582000
rect 154000 580000 245900 581400
rect 283800 580600 285400 594000
rect 286000 580600 287600 602000
rect -800 564220 1660 564242
rect -800 564057 4430 564220
rect -800 559593 888 564057
rect 4232 559593 4430 564057
rect -800 559442 4430 559593
rect 680 554972 4430 559442
rect 680 554242 1028 554972
rect -800 550028 1028 554242
rect 3972 550028 4430 554972
rect -800 549442 4430 550028
rect 680 549410 4430 549442
rect 260 508118 57120 508140
rect 260 508096 57022 508118
rect -800 508062 57022 508096
rect 57078 508062 57120 508118
rect -800 508038 57120 508062
rect -800 507984 57022 508038
rect 260 507982 57022 507984
rect 57078 507982 57120 508038
rect 260 507960 57120 507982
rect 280 466078 56860 466100
rect 280 466056 56762 466078
rect -800 466022 56762 466056
rect 56818 466022 56860 466078
rect -800 465998 56860 466022
rect -800 465944 56762 465998
rect 280 465942 56762 465944
rect 56818 465942 56860 465998
rect 280 465920 56860 465942
rect 360 421658 56620 421680
rect 360 421652 56522 421658
rect -800 421602 56522 421652
rect 56578 421602 56620 421658
rect -800 421578 56620 421602
rect -800 421540 56522 421578
rect 360 421522 56522 421540
rect 56578 421522 56620 421578
rect 360 421500 56620 421522
rect 400 378458 56340 378480
rect 400 378430 56242 378458
rect -800 378402 56242 378430
rect 56298 378402 56340 378458
rect -800 378378 56340 378402
rect -800 378322 56242 378378
rect 56298 378322 56340 378378
rect -800 378318 56340 378322
rect 400 378300 56340 378318
rect 260 335218 56100 335240
rect 260 335208 56002 335218
rect -800 335162 56002 335208
rect 56058 335162 56100 335218
rect -800 335138 56100 335162
rect -800 335096 56002 335138
rect 260 335082 56002 335096
rect 56058 335082 56100 335138
rect 260 335060 56100 335082
rect 200 295532 800 295600
rect -800 295420 800 295532
rect 200 295400 800 295420
rect 154000 295400 158000 580000
rect 200 294600 158000 295400
rect 200 294350 800 294600
rect -800 294238 800 294350
rect 200 294200 800 294238
rect 154000 294000 158000 294600
rect 1650 177690 20600 178000
rect 982 177688 20600 177690
rect -800 177582 20600 177688
rect -800 172888 11628 177582
rect 982 172318 11628 172888
rect 20172 172318 20600 177582
rect 982 171900 20600 172318
rect 982 167688 5298 171900
rect -800 162890 5298 167688
rect -800 162888 1660 162890
<< via3 >>
rect 42598 688413 43142 689437
rect 40773 676133 41637 677237
rect 23218 668688 23362 669072
rect 73008 635008 78992 646992
rect 173628 699628 175372 701772
rect 511008 694008 524992 701992
rect 572008 631008 579992 642992
rect 22008 604008 23992 605992
rect 165028 583028 181972 589972
rect 888 559593 4232 564057
rect 1028 550028 3972 554972
rect 11628 172318 20172 177582
<< metal4 >>
rect 165594 703000 170594 704800
rect 175894 703000 180894 704800
rect 165000 701772 182000 703000
rect 165000 699628 173628 701772
rect 175372 699628 182000 701772
rect 42500 689437 43450 689470
rect 42500 688413 42598 689437
rect 43142 688413 43450 689437
rect 42500 677320 43450 688413
rect 40720 677237 43450 677320
rect 40720 676133 40773 677237
rect 41637 676133 43450 677237
rect 40720 676090 43450 676133
rect 40720 676080 43220 676090
rect 60220 676010 65450 676030
rect 56870 675823 65450 676010
rect 56870 675587 60947 675823
rect 61183 675587 61267 675823
rect 61503 675587 61587 675823
rect 61823 675587 61907 675823
rect 62143 675587 62227 675823
rect 62463 675587 62547 675823
rect 62783 675587 62867 675823
rect 63103 675587 63187 675823
rect 63423 675587 63507 675823
rect 63743 675587 63827 675823
rect 64063 675587 64147 675823
rect 64383 675587 64467 675823
rect 64703 675587 64787 675823
rect 65023 675587 65107 675823
rect 65343 675587 65450 675823
rect 56870 675370 65450 675587
rect 23190 669072 23390 669110
rect 23190 668688 23218 669072
rect 23362 668688 23390 669072
rect 23190 608120 23390 668688
rect 26600 633690 28120 662640
rect 72999 646992 79001 647001
rect 72999 646878 73008 646992
rect 78992 646878 79001 646992
rect 72999 635122 73002 646878
rect 78998 635122 79001 646878
rect 72999 635008 73008 635122
rect 78992 635008 79001 635122
rect 72999 634999 79001 635008
rect 26090 633478 28790 633690
rect 26090 631642 26347 633478
rect 28503 631642 28790 633478
rect 26090 631490 28790 631642
rect 32100 620173 39650 620900
rect 32100 614177 32937 620173
rect 38613 614177 39650 620173
rect 32100 613600 39650 614177
rect 21660 605992 25780 608120
rect 21660 604008 22008 605992
rect 23992 604008 25780 605992
rect 21660 603350 25780 604008
rect 690 564057 4450 564270
rect 690 559593 888 564057
rect 4232 559593 4450 564057
rect 690 559400 4450 559593
rect 999 554972 4001 555001
rect 999 550028 1028 554972
rect 3972 550028 4001 554972
rect 999 549999 4001 550028
rect 30150 178000 39650 613600
rect 165000 590001 182000 699628
rect 510000 701992 526000 703000
rect 510000 694008 511008 701992
rect 524992 694008 526000 701992
rect 305500 644958 316500 646500
rect 238000 643958 248000 644000
rect 238000 636042 238082 643958
rect 247918 636042 248000 643958
rect 164999 589972 182001 590001
rect 164999 583028 165028 589972
rect 181972 583028 182001 589972
rect 164999 582999 182001 583028
rect 238000 584000 248000 636042
rect 305500 637042 307042 644958
rect 314958 637042 316500 644958
rect 238000 580000 260000 584000
rect 305500 580300 316500 637042
rect 238200 570900 240100 574000
rect 258800 571400 260000 580000
rect 238200 568100 239300 570900
rect 238200 563688 240200 568100
rect 238200 558012 238352 563688
rect 239548 558012 240200 563688
rect 510000 562958 526000 694008
rect 570000 642992 582000 645000
rect 570000 631008 572008 642992
rect 579992 631008 582000 642992
rect 570000 630000 582000 631008
rect 238200 558000 240200 558012
rect 263600 557748 316600 558100
rect 263600 556552 263742 557748
rect 316458 556552 316600 557748
rect 263600 556400 316600 556552
rect 510000 555042 511002 562958
rect 524998 555042 526000 562958
rect 510000 554000 526000 555042
rect 11100 177582 39650 178000
rect 11100 172318 11628 177582
rect 20172 172318 39650 177582
rect 11100 171950 39650 172318
rect 11100 171900 34150 171950
<< via4 >>
rect 60947 675587 61183 675823
rect 61267 675587 61503 675823
rect 61587 675587 61823 675823
rect 61907 675587 62143 675823
rect 62227 675587 62463 675823
rect 62547 675587 62783 675823
rect 62867 675587 63103 675823
rect 63187 675587 63423 675823
rect 63507 675587 63743 675823
rect 63827 675587 64063 675823
rect 64147 675587 64383 675823
rect 64467 675587 64703 675823
rect 64787 675587 65023 675823
rect 65107 675587 65343 675823
rect 73002 635122 73008 646878
rect 73008 635122 78992 646878
rect 78992 635122 78998 646878
rect 26347 631642 28503 633478
rect 32937 614177 38613 620173
rect 1002 559627 4118 564023
rect 1102 550142 3898 554858
rect 238082 636042 247918 643958
rect 307042 637042 314958 644958
rect 238352 558012 239548 563688
rect 572042 631122 579958 642878
rect 263742 556552 316458 557748
rect 511002 555042 524998 562958
<< metal5 >>
rect 165594 702300 170594 704800
rect 175894 702300 180894 704800
rect 60790 675823 65590 676060
rect 60790 675587 60947 675823
rect 61183 675587 61267 675823
rect 61503 675587 61587 675823
rect 61823 675587 61907 675823
rect 62143 675587 62227 675823
rect 62463 675587 62547 675823
rect 62783 675587 62867 675823
rect 63103 675587 63187 675823
rect 63423 675587 63507 675823
rect 63743 675587 63827 675823
rect 64063 675587 64147 675823
rect 64383 675587 64467 675823
rect 64703 675587 64787 675823
rect 65023 675587 65107 675823
rect 65343 675587 65590 675823
rect 26080 633478 28810 633710
rect 26080 631642 26347 633478
rect 28503 631642 28810 633478
rect 26080 564330 28810 631642
rect 33890 625850 34330 675040
rect 39240 625850 39680 674940
rect 42370 625850 42840 674830
rect 44740 625850 45180 675000
rect 45790 625850 46240 663160
rect 60790 652300 65590 675587
rect 32150 620173 51000 625850
rect 32150 614177 32937 620173
rect 38613 614177 51000 620173
rect 32150 613550 51000 614177
rect 60820 564330 65590 652300
rect 72976 647000 79024 647024
rect 72976 646878 582000 647000
rect 72976 635122 73002 646878
rect 78998 644958 582000 646878
rect 78998 643958 307042 644958
rect 78998 636042 238082 643958
rect 247918 637042 307042 643958
rect 314958 642878 582000 644958
rect 314958 637042 572042 642878
rect 247918 636042 572042 637042
rect 78998 635122 572042 636042
rect 72976 635000 572042 635122
rect 72976 634976 79024 635000
rect 564000 631122 572042 635000
rect 579958 631122 582000 642878
rect 564000 630000 582000 631122
rect 26080 564320 65590 564330
rect 1770 564270 65590 564320
rect 690 564023 65590 564270
rect 690 559627 1002 564023
rect 4118 564000 65590 564023
rect 4118 563688 526000 564000
rect 4118 559627 238352 563688
rect 690 559400 238352 559627
rect 1000 558012 238352 559400
rect 239548 562958 526000 563688
rect 239548 558012 511002 562958
rect 1000 557748 511002 558012
rect 1000 556552 263742 557748
rect 316458 556552 511002 557748
rect 1000 555042 511002 556552
rect 524998 555042 526000 562958
rect 1000 555024 526000 555042
rect 976 554858 526000 555024
rect 976 550142 1102 554858
rect 3898 550142 526000 554858
rect 976 550000 526000 550142
rect 976 549976 4024 550000
use BGR_lvs  BGR_lvs_0
timestamp 1663011646
transform 1 0 254230 0 1 568403
box -14220 -10400 62400 12600
use VCO  VCO_0
timestamp 1663011646
transform 1 0 -7837 0 1 638742
box 31151 20430 65400 41670
<< labels >>
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1400 0 0 0 io_analog[10]
port 1 nsew
flabel metal5 s 26080 559400 65590 564330 0 FreeSans 20000 0 0 0 GND
port 2 nsew
rlabel metal2 s 56980 508120 57120 660100 4 CTRL1
port 3 nsew
rlabel metal2 s 56720 466080 56860 660460 4 CTRL2
port 4 nsew
rlabel metal2 s 56480 421660 56620 660980 4 CTRL3
port 5 nsew
rlabel metal2 s 56200 378460 56340 661580 4 CTRL4
port 6 nsew
rlabel metal2 s 55960 335220 56100 662500 4 CTRL5
port 7 nsew
flabel metal1 s 14920 668060 15420 682040 0 FreeSans 10000 0 0 0 VCTRL
port 8 nsew
flabel metal4 s 21660 603350 25780 608120 0 FreeSans 10000 0 0 0 REF
port 9 nsew
rlabel metal3 s 17070 688210 41870 689330 4 OUT0
port 10 nsew
rlabel metal3 s 43180 688360 70760 689480 4 OUT180
port 11 nsew
flabel metal3 s -800 295420 480 295532 0 FreeSans 1400 0 0 0 gpio_analog[12]
port 12 nsew
flabel metal3 s -800 294238 480 294350 0 FreeSans 1400 0 0 0 gpio_noesd[12]
port 13 nsew
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal4 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal5 s 175894 702300 180894 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 2400 180 0 0 io_analog[7]
port 15 nsew
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 2400 180 0 0 io_analog[8]
port 16 nsew
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 2400 180 0 0 io_analog[9]
port 17 nsew
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal4 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal5 s 165594 702300 170594 704800 0 FreeSans 2400 180 0 0 io_analog[6]
port 14 nsew
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 2400 180 0 0 io_clamp_high[2]
port 18 nsew
flabel metal3 s -800 507984 480 508096 0 FreeSans 1400 0 0 0 io_in[14]
port 19 nsew
flabel metal3 s -800 421540 480 421652 0 FreeSans 1400 0 0 0 io_in[16]
port 20 nsew
flabel metal3 s -800 378318 480 378430 0 FreeSans 1400 0 0 0 io_in[17]
port 21 nsew
flabel metal3 s -800 335096 480 335208 0 FreeSans 1400 0 0 0 io_in[18]
port 22 nsew
flabel metal3 s -800 465944 480 466056 0 FreeSans 1400 0 0 0 io_in_3v3[15]
port 23 nsew
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1400 0 0 0 vccd1
port 24 nsew
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1400 0 0 0 vccd1
port 24 nsew
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1400 0 0 0 vccd2
port 25 nsew
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1400 0 0 0 vccd2
port 25 nsew
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 2400 180 0 0 vssa1
port 26 nsew
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 2400 180 0 0 vssa1
port 26 nsew
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1400 0 0 0 vssa2
port 27 nsew
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1400 0 0 0 vssa2
port 27 nsew
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1400 0 0 0 vssd2
port 28 nsew
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1400 0 0 0 vssd2
port 28 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
