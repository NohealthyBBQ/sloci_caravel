magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -812 -284 812 284
<< pmoslvt >>
rect -616 -64 -416 136
rect -358 -64 -158 136
rect -100 -64 100 136
rect 158 -64 358 136
rect 416 -64 616 136
<< pdiff >>
rect -674 121 -616 136
rect -674 87 -662 121
rect -628 87 -616 121
rect -674 53 -616 87
rect -674 19 -662 53
rect -628 19 -616 53
rect -674 -15 -616 19
rect -674 -49 -662 -15
rect -628 -49 -616 -15
rect -674 -64 -616 -49
rect -416 121 -358 136
rect -416 87 -404 121
rect -370 87 -358 121
rect -416 53 -358 87
rect -416 19 -404 53
rect -370 19 -358 53
rect -416 -15 -358 19
rect -416 -49 -404 -15
rect -370 -49 -358 -15
rect -416 -64 -358 -49
rect -158 121 -100 136
rect -158 87 -146 121
rect -112 87 -100 121
rect -158 53 -100 87
rect -158 19 -146 53
rect -112 19 -100 53
rect -158 -15 -100 19
rect -158 -49 -146 -15
rect -112 -49 -100 -15
rect -158 -64 -100 -49
rect 100 121 158 136
rect 100 87 112 121
rect 146 87 158 121
rect 100 53 158 87
rect 100 19 112 53
rect 146 19 158 53
rect 100 -15 158 19
rect 100 -49 112 -15
rect 146 -49 158 -15
rect 100 -64 158 -49
rect 358 121 416 136
rect 358 87 370 121
rect 404 87 416 121
rect 358 53 416 87
rect 358 19 370 53
rect 404 19 416 53
rect 358 -15 416 19
rect 358 -49 370 -15
rect 404 -49 416 -15
rect 358 -64 416 -49
rect 616 121 674 136
rect 616 87 628 121
rect 662 87 674 121
rect 616 53 674 87
rect 616 19 628 53
rect 662 19 674 53
rect 616 -15 674 19
rect 616 -49 628 -15
rect 662 -49 674 -15
rect 616 -64 674 -49
<< pdiffc >>
rect -662 87 -628 121
rect -662 19 -628 53
rect -662 -49 -628 -15
rect -404 87 -370 121
rect -404 19 -370 53
rect -404 -49 -370 -15
rect -146 87 -112 121
rect -146 19 -112 53
rect -146 -49 -112 -15
rect 112 87 146 121
rect 112 19 146 53
rect 112 -49 146 -15
rect 370 87 404 121
rect 370 19 404 53
rect 370 -49 404 -15
rect 628 87 662 121
rect 628 19 662 53
rect 628 -49 662 -15
<< nsubdiff >>
rect -776 214 776 248
rect -776 119 -742 214
rect -776 51 -742 85
rect -776 -17 -742 17
rect -776 -85 -742 -51
rect 742 119 776 214
rect 742 51 776 85
rect 742 -17 776 17
rect -776 -214 -742 -119
rect 742 -85 776 -51
rect 742 -214 776 -119
rect -776 -248 776 -214
<< nsubdiffcont >>
rect -776 85 -742 119
rect -776 17 -742 51
rect -776 -51 -742 -17
rect 742 85 776 119
rect 742 17 776 51
rect 742 -51 776 -17
rect -776 -119 -742 -85
rect 742 -119 776 -85
<< poly >>
rect -616 136 -416 162
rect -358 136 -158 162
rect -100 136 100 162
rect 158 136 358 162
rect 416 136 616 162
rect -616 -111 -416 -64
rect -616 -145 -567 -111
rect -533 -145 -499 -111
rect -465 -145 -416 -111
rect -616 -161 -416 -145
rect -358 -111 -158 -64
rect -358 -145 -309 -111
rect -275 -145 -241 -111
rect -207 -145 -158 -111
rect -358 -161 -158 -145
rect -100 -111 100 -64
rect -100 -145 -51 -111
rect -17 -145 17 -111
rect 51 -145 100 -111
rect -100 -161 100 -145
rect 158 -111 358 -64
rect 158 -145 207 -111
rect 241 -145 275 -111
rect 309 -145 358 -111
rect 158 -161 358 -145
rect 416 -111 616 -64
rect 416 -145 465 -111
rect 499 -145 533 -111
rect 567 -145 616 -111
rect 416 -161 616 -145
<< polycont >>
rect -567 -145 -533 -111
rect -499 -145 -465 -111
rect -309 -145 -275 -111
rect -241 -145 -207 -111
rect -51 -145 -17 -111
rect 17 -145 51 -111
rect 207 -145 241 -111
rect 275 -145 309 -111
rect 465 -145 499 -111
rect 533 -145 567 -111
<< locali >>
rect -776 214 776 248
rect -776 119 -742 214
rect -776 51 -742 85
rect -776 -17 -742 17
rect -776 -85 -742 -51
rect -662 121 -628 140
rect -662 53 -628 55
rect -662 17 -628 19
rect -662 -68 -628 -49
rect -404 121 -370 140
rect -404 53 -370 55
rect -404 17 -370 19
rect -404 -68 -370 -49
rect -146 121 -112 140
rect -146 53 -112 55
rect -146 17 -112 19
rect -146 -68 -112 -49
rect 112 121 146 140
rect 112 53 146 55
rect 112 17 146 19
rect 112 -68 146 -49
rect 370 121 404 140
rect 370 53 404 55
rect 370 17 404 19
rect 370 -68 404 -49
rect 628 121 662 140
rect 628 53 662 55
rect 628 17 662 19
rect 628 -68 662 -49
rect 742 119 776 214
rect 742 51 776 85
rect 742 -17 776 17
rect 742 -85 776 -51
rect -776 -214 -742 -119
rect -616 -145 -569 -111
rect -533 -145 -499 -111
rect -463 -145 -416 -111
rect -358 -145 -311 -111
rect -275 -145 -241 -111
rect -205 -145 -158 -111
rect -100 -145 -53 -111
rect -17 -145 17 -111
rect 53 -145 100 -111
rect 158 -145 205 -111
rect 241 -145 275 -111
rect 311 -145 358 -111
rect 416 -145 463 -111
rect 499 -145 533 -111
rect 569 -145 616 -111
rect 742 -214 776 -119
rect -776 -248 776 -214
<< viali >>
rect -662 87 -628 89
rect -662 55 -628 87
rect -662 -15 -628 17
rect -662 -17 -628 -15
rect -404 87 -370 89
rect -404 55 -370 87
rect -404 -15 -370 17
rect -404 -17 -370 -15
rect -146 87 -112 89
rect -146 55 -112 87
rect -146 -15 -112 17
rect -146 -17 -112 -15
rect 112 87 146 89
rect 112 55 146 87
rect 112 -15 146 17
rect 112 -17 146 -15
rect 370 87 404 89
rect 370 55 404 87
rect 370 -15 404 17
rect 370 -17 404 -15
rect 628 87 662 89
rect 628 55 662 87
rect 628 -15 662 17
rect 628 -17 662 -15
rect -569 -145 -567 -111
rect -567 -145 -535 -111
rect -497 -145 -465 -111
rect -465 -145 -463 -111
rect -311 -145 -309 -111
rect -309 -145 -277 -111
rect -239 -145 -207 -111
rect -207 -145 -205 -111
rect -53 -145 -51 -111
rect -51 -145 -19 -111
rect 19 -145 51 -111
rect 51 -145 53 -111
rect 205 -145 207 -111
rect 207 -145 239 -111
rect 277 -145 309 -111
rect 309 -145 311 -111
rect 463 -145 465 -111
rect 465 -145 497 -111
rect 535 -145 567 -111
rect 567 -145 569 -111
<< metal1 >>
rect -668 89 -622 136
rect -668 55 -662 89
rect -628 55 -622 89
rect -668 17 -622 55
rect -668 -17 -662 17
rect -628 -17 -622 17
rect -668 -64 -622 -17
rect -410 89 -364 136
rect -410 55 -404 89
rect -370 55 -364 89
rect -410 17 -364 55
rect -410 -17 -404 17
rect -370 -17 -364 17
rect -410 -64 -364 -17
rect -152 89 -106 136
rect -152 55 -146 89
rect -112 55 -106 89
rect -152 17 -106 55
rect -152 -17 -146 17
rect -112 -17 -106 17
rect -152 -64 -106 -17
rect 106 89 152 136
rect 106 55 112 89
rect 146 55 152 89
rect 106 17 152 55
rect 106 -17 112 17
rect 146 -17 152 17
rect 106 -64 152 -17
rect 364 89 410 136
rect 364 55 370 89
rect 404 55 410 89
rect 364 17 410 55
rect 364 -17 370 17
rect 404 -17 410 17
rect 364 -64 410 -17
rect 622 89 668 136
rect 622 55 628 89
rect 662 55 668 89
rect 622 17 668 55
rect 622 -17 628 17
rect 662 -17 668 17
rect 622 -64 668 -17
rect -612 -111 -420 -105
rect -612 -145 -569 -111
rect -535 -145 -497 -111
rect -463 -145 -420 -111
rect -612 -151 -420 -145
rect -354 -111 -162 -105
rect -354 -145 -311 -111
rect -277 -145 -239 -111
rect -205 -145 -162 -111
rect -354 -151 -162 -145
rect -96 -111 96 -105
rect -96 -145 -53 -111
rect -19 -145 19 -111
rect 53 -145 96 -111
rect -96 -151 96 -145
rect 162 -111 354 -105
rect 162 -145 205 -111
rect 239 -145 277 -111
rect 311 -145 354 -111
rect 162 -151 354 -145
rect 420 -111 612 -105
rect 420 -145 463 -111
rect 497 -145 535 -111
rect 569 -145 612 -111
rect 420 -151 612 -145
<< properties >>
string FIXED_BBOX -759 -231 759 231
<< end >>
