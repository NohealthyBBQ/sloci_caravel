magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -1273 -2831 1273 2831
<< pmoslvt >>
rect -1077 1483 -977 2683
rect -919 1483 -819 2683
rect -761 1483 -661 2683
rect -603 1483 -503 2683
rect -445 1483 -345 2683
rect -287 1483 -187 2683
rect -129 1483 -29 2683
rect 29 1483 129 2683
rect 187 1483 287 2683
rect 345 1483 445 2683
rect 503 1483 603 2683
rect 661 1483 761 2683
rect 819 1483 919 2683
rect 977 1483 1077 2683
rect -1077 118 -977 1318
rect -919 118 -819 1318
rect -761 118 -661 1318
rect -603 118 -503 1318
rect -445 118 -345 1318
rect -287 118 -187 1318
rect -129 118 -29 1318
rect 29 118 129 1318
rect 187 118 287 1318
rect 345 118 445 1318
rect 503 118 603 1318
rect 661 118 761 1318
rect 819 118 919 1318
rect 977 118 1077 1318
rect -1077 -1247 -977 -47
rect -919 -1247 -819 -47
rect -761 -1247 -661 -47
rect -603 -1247 -503 -47
rect -445 -1247 -345 -47
rect -287 -1247 -187 -47
rect -129 -1247 -29 -47
rect 29 -1247 129 -47
rect 187 -1247 287 -47
rect 345 -1247 445 -47
rect 503 -1247 603 -47
rect 661 -1247 761 -47
rect 819 -1247 919 -47
rect 977 -1247 1077 -47
rect -1077 -2612 -977 -1412
rect -919 -2612 -819 -1412
rect -761 -2612 -661 -1412
rect -603 -2612 -503 -1412
rect -445 -2612 -345 -1412
rect -287 -2612 -187 -1412
rect -129 -2612 -29 -1412
rect 29 -2612 129 -1412
rect 187 -2612 287 -1412
rect 345 -2612 445 -1412
rect 503 -2612 603 -1412
rect 661 -2612 761 -1412
rect 819 -2612 919 -1412
rect 977 -2612 1077 -1412
<< pdiff >>
rect -1135 2644 -1077 2683
rect -1135 2610 -1123 2644
rect -1089 2610 -1077 2644
rect -1135 2576 -1077 2610
rect -1135 2542 -1123 2576
rect -1089 2542 -1077 2576
rect -1135 2508 -1077 2542
rect -1135 2474 -1123 2508
rect -1089 2474 -1077 2508
rect -1135 2440 -1077 2474
rect -1135 2406 -1123 2440
rect -1089 2406 -1077 2440
rect -1135 2372 -1077 2406
rect -1135 2338 -1123 2372
rect -1089 2338 -1077 2372
rect -1135 2304 -1077 2338
rect -1135 2270 -1123 2304
rect -1089 2270 -1077 2304
rect -1135 2236 -1077 2270
rect -1135 2202 -1123 2236
rect -1089 2202 -1077 2236
rect -1135 2168 -1077 2202
rect -1135 2134 -1123 2168
rect -1089 2134 -1077 2168
rect -1135 2100 -1077 2134
rect -1135 2066 -1123 2100
rect -1089 2066 -1077 2100
rect -1135 2032 -1077 2066
rect -1135 1998 -1123 2032
rect -1089 1998 -1077 2032
rect -1135 1964 -1077 1998
rect -1135 1930 -1123 1964
rect -1089 1930 -1077 1964
rect -1135 1896 -1077 1930
rect -1135 1862 -1123 1896
rect -1089 1862 -1077 1896
rect -1135 1828 -1077 1862
rect -1135 1794 -1123 1828
rect -1089 1794 -1077 1828
rect -1135 1760 -1077 1794
rect -1135 1726 -1123 1760
rect -1089 1726 -1077 1760
rect -1135 1692 -1077 1726
rect -1135 1658 -1123 1692
rect -1089 1658 -1077 1692
rect -1135 1624 -1077 1658
rect -1135 1590 -1123 1624
rect -1089 1590 -1077 1624
rect -1135 1556 -1077 1590
rect -1135 1522 -1123 1556
rect -1089 1522 -1077 1556
rect -1135 1483 -1077 1522
rect -977 2644 -919 2683
rect -977 2610 -965 2644
rect -931 2610 -919 2644
rect -977 2576 -919 2610
rect -977 2542 -965 2576
rect -931 2542 -919 2576
rect -977 2508 -919 2542
rect -977 2474 -965 2508
rect -931 2474 -919 2508
rect -977 2440 -919 2474
rect -977 2406 -965 2440
rect -931 2406 -919 2440
rect -977 2372 -919 2406
rect -977 2338 -965 2372
rect -931 2338 -919 2372
rect -977 2304 -919 2338
rect -977 2270 -965 2304
rect -931 2270 -919 2304
rect -977 2236 -919 2270
rect -977 2202 -965 2236
rect -931 2202 -919 2236
rect -977 2168 -919 2202
rect -977 2134 -965 2168
rect -931 2134 -919 2168
rect -977 2100 -919 2134
rect -977 2066 -965 2100
rect -931 2066 -919 2100
rect -977 2032 -919 2066
rect -977 1998 -965 2032
rect -931 1998 -919 2032
rect -977 1964 -919 1998
rect -977 1930 -965 1964
rect -931 1930 -919 1964
rect -977 1896 -919 1930
rect -977 1862 -965 1896
rect -931 1862 -919 1896
rect -977 1828 -919 1862
rect -977 1794 -965 1828
rect -931 1794 -919 1828
rect -977 1760 -919 1794
rect -977 1726 -965 1760
rect -931 1726 -919 1760
rect -977 1692 -919 1726
rect -977 1658 -965 1692
rect -931 1658 -919 1692
rect -977 1624 -919 1658
rect -977 1590 -965 1624
rect -931 1590 -919 1624
rect -977 1556 -919 1590
rect -977 1522 -965 1556
rect -931 1522 -919 1556
rect -977 1483 -919 1522
rect -819 2644 -761 2683
rect -819 2610 -807 2644
rect -773 2610 -761 2644
rect -819 2576 -761 2610
rect -819 2542 -807 2576
rect -773 2542 -761 2576
rect -819 2508 -761 2542
rect -819 2474 -807 2508
rect -773 2474 -761 2508
rect -819 2440 -761 2474
rect -819 2406 -807 2440
rect -773 2406 -761 2440
rect -819 2372 -761 2406
rect -819 2338 -807 2372
rect -773 2338 -761 2372
rect -819 2304 -761 2338
rect -819 2270 -807 2304
rect -773 2270 -761 2304
rect -819 2236 -761 2270
rect -819 2202 -807 2236
rect -773 2202 -761 2236
rect -819 2168 -761 2202
rect -819 2134 -807 2168
rect -773 2134 -761 2168
rect -819 2100 -761 2134
rect -819 2066 -807 2100
rect -773 2066 -761 2100
rect -819 2032 -761 2066
rect -819 1998 -807 2032
rect -773 1998 -761 2032
rect -819 1964 -761 1998
rect -819 1930 -807 1964
rect -773 1930 -761 1964
rect -819 1896 -761 1930
rect -819 1862 -807 1896
rect -773 1862 -761 1896
rect -819 1828 -761 1862
rect -819 1794 -807 1828
rect -773 1794 -761 1828
rect -819 1760 -761 1794
rect -819 1726 -807 1760
rect -773 1726 -761 1760
rect -819 1692 -761 1726
rect -819 1658 -807 1692
rect -773 1658 -761 1692
rect -819 1624 -761 1658
rect -819 1590 -807 1624
rect -773 1590 -761 1624
rect -819 1556 -761 1590
rect -819 1522 -807 1556
rect -773 1522 -761 1556
rect -819 1483 -761 1522
rect -661 2644 -603 2683
rect -661 2610 -649 2644
rect -615 2610 -603 2644
rect -661 2576 -603 2610
rect -661 2542 -649 2576
rect -615 2542 -603 2576
rect -661 2508 -603 2542
rect -661 2474 -649 2508
rect -615 2474 -603 2508
rect -661 2440 -603 2474
rect -661 2406 -649 2440
rect -615 2406 -603 2440
rect -661 2372 -603 2406
rect -661 2338 -649 2372
rect -615 2338 -603 2372
rect -661 2304 -603 2338
rect -661 2270 -649 2304
rect -615 2270 -603 2304
rect -661 2236 -603 2270
rect -661 2202 -649 2236
rect -615 2202 -603 2236
rect -661 2168 -603 2202
rect -661 2134 -649 2168
rect -615 2134 -603 2168
rect -661 2100 -603 2134
rect -661 2066 -649 2100
rect -615 2066 -603 2100
rect -661 2032 -603 2066
rect -661 1998 -649 2032
rect -615 1998 -603 2032
rect -661 1964 -603 1998
rect -661 1930 -649 1964
rect -615 1930 -603 1964
rect -661 1896 -603 1930
rect -661 1862 -649 1896
rect -615 1862 -603 1896
rect -661 1828 -603 1862
rect -661 1794 -649 1828
rect -615 1794 -603 1828
rect -661 1760 -603 1794
rect -661 1726 -649 1760
rect -615 1726 -603 1760
rect -661 1692 -603 1726
rect -661 1658 -649 1692
rect -615 1658 -603 1692
rect -661 1624 -603 1658
rect -661 1590 -649 1624
rect -615 1590 -603 1624
rect -661 1556 -603 1590
rect -661 1522 -649 1556
rect -615 1522 -603 1556
rect -661 1483 -603 1522
rect -503 2644 -445 2683
rect -503 2610 -491 2644
rect -457 2610 -445 2644
rect -503 2576 -445 2610
rect -503 2542 -491 2576
rect -457 2542 -445 2576
rect -503 2508 -445 2542
rect -503 2474 -491 2508
rect -457 2474 -445 2508
rect -503 2440 -445 2474
rect -503 2406 -491 2440
rect -457 2406 -445 2440
rect -503 2372 -445 2406
rect -503 2338 -491 2372
rect -457 2338 -445 2372
rect -503 2304 -445 2338
rect -503 2270 -491 2304
rect -457 2270 -445 2304
rect -503 2236 -445 2270
rect -503 2202 -491 2236
rect -457 2202 -445 2236
rect -503 2168 -445 2202
rect -503 2134 -491 2168
rect -457 2134 -445 2168
rect -503 2100 -445 2134
rect -503 2066 -491 2100
rect -457 2066 -445 2100
rect -503 2032 -445 2066
rect -503 1998 -491 2032
rect -457 1998 -445 2032
rect -503 1964 -445 1998
rect -503 1930 -491 1964
rect -457 1930 -445 1964
rect -503 1896 -445 1930
rect -503 1862 -491 1896
rect -457 1862 -445 1896
rect -503 1828 -445 1862
rect -503 1794 -491 1828
rect -457 1794 -445 1828
rect -503 1760 -445 1794
rect -503 1726 -491 1760
rect -457 1726 -445 1760
rect -503 1692 -445 1726
rect -503 1658 -491 1692
rect -457 1658 -445 1692
rect -503 1624 -445 1658
rect -503 1590 -491 1624
rect -457 1590 -445 1624
rect -503 1556 -445 1590
rect -503 1522 -491 1556
rect -457 1522 -445 1556
rect -503 1483 -445 1522
rect -345 2644 -287 2683
rect -345 2610 -333 2644
rect -299 2610 -287 2644
rect -345 2576 -287 2610
rect -345 2542 -333 2576
rect -299 2542 -287 2576
rect -345 2508 -287 2542
rect -345 2474 -333 2508
rect -299 2474 -287 2508
rect -345 2440 -287 2474
rect -345 2406 -333 2440
rect -299 2406 -287 2440
rect -345 2372 -287 2406
rect -345 2338 -333 2372
rect -299 2338 -287 2372
rect -345 2304 -287 2338
rect -345 2270 -333 2304
rect -299 2270 -287 2304
rect -345 2236 -287 2270
rect -345 2202 -333 2236
rect -299 2202 -287 2236
rect -345 2168 -287 2202
rect -345 2134 -333 2168
rect -299 2134 -287 2168
rect -345 2100 -287 2134
rect -345 2066 -333 2100
rect -299 2066 -287 2100
rect -345 2032 -287 2066
rect -345 1998 -333 2032
rect -299 1998 -287 2032
rect -345 1964 -287 1998
rect -345 1930 -333 1964
rect -299 1930 -287 1964
rect -345 1896 -287 1930
rect -345 1862 -333 1896
rect -299 1862 -287 1896
rect -345 1828 -287 1862
rect -345 1794 -333 1828
rect -299 1794 -287 1828
rect -345 1760 -287 1794
rect -345 1726 -333 1760
rect -299 1726 -287 1760
rect -345 1692 -287 1726
rect -345 1658 -333 1692
rect -299 1658 -287 1692
rect -345 1624 -287 1658
rect -345 1590 -333 1624
rect -299 1590 -287 1624
rect -345 1556 -287 1590
rect -345 1522 -333 1556
rect -299 1522 -287 1556
rect -345 1483 -287 1522
rect -187 2644 -129 2683
rect -187 2610 -175 2644
rect -141 2610 -129 2644
rect -187 2576 -129 2610
rect -187 2542 -175 2576
rect -141 2542 -129 2576
rect -187 2508 -129 2542
rect -187 2474 -175 2508
rect -141 2474 -129 2508
rect -187 2440 -129 2474
rect -187 2406 -175 2440
rect -141 2406 -129 2440
rect -187 2372 -129 2406
rect -187 2338 -175 2372
rect -141 2338 -129 2372
rect -187 2304 -129 2338
rect -187 2270 -175 2304
rect -141 2270 -129 2304
rect -187 2236 -129 2270
rect -187 2202 -175 2236
rect -141 2202 -129 2236
rect -187 2168 -129 2202
rect -187 2134 -175 2168
rect -141 2134 -129 2168
rect -187 2100 -129 2134
rect -187 2066 -175 2100
rect -141 2066 -129 2100
rect -187 2032 -129 2066
rect -187 1998 -175 2032
rect -141 1998 -129 2032
rect -187 1964 -129 1998
rect -187 1930 -175 1964
rect -141 1930 -129 1964
rect -187 1896 -129 1930
rect -187 1862 -175 1896
rect -141 1862 -129 1896
rect -187 1828 -129 1862
rect -187 1794 -175 1828
rect -141 1794 -129 1828
rect -187 1760 -129 1794
rect -187 1726 -175 1760
rect -141 1726 -129 1760
rect -187 1692 -129 1726
rect -187 1658 -175 1692
rect -141 1658 -129 1692
rect -187 1624 -129 1658
rect -187 1590 -175 1624
rect -141 1590 -129 1624
rect -187 1556 -129 1590
rect -187 1522 -175 1556
rect -141 1522 -129 1556
rect -187 1483 -129 1522
rect -29 2644 29 2683
rect -29 2610 -17 2644
rect 17 2610 29 2644
rect -29 2576 29 2610
rect -29 2542 -17 2576
rect 17 2542 29 2576
rect -29 2508 29 2542
rect -29 2474 -17 2508
rect 17 2474 29 2508
rect -29 2440 29 2474
rect -29 2406 -17 2440
rect 17 2406 29 2440
rect -29 2372 29 2406
rect -29 2338 -17 2372
rect 17 2338 29 2372
rect -29 2304 29 2338
rect -29 2270 -17 2304
rect 17 2270 29 2304
rect -29 2236 29 2270
rect -29 2202 -17 2236
rect 17 2202 29 2236
rect -29 2168 29 2202
rect -29 2134 -17 2168
rect 17 2134 29 2168
rect -29 2100 29 2134
rect -29 2066 -17 2100
rect 17 2066 29 2100
rect -29 2032 29 2066
rect -29 1998 -17 2032
rect 17 1998 29 2032
rect -29 1964 29 1998
rect -29 1930 -17 1964
rect 17 1930 29 1964
rect -29 1896 29 1930
rect -29 1862 -17 1896
rect 17 1862 29 1896
rect -29 1828 29 1862
rect -29 1794 -17 1828
rect 17 1794 29 1828
rect -29 1760 29 1794
rect -29 1726 -17 1760
rect 17 1726 29 1760
rect -29 1692 29 1726
rect -29 1658 -17 1692
rect 17 1658 29 1692
rect -29 1624 29 1658
rect -29 1590 -17 1624
rect 17 1590 29 1624
rect -29 1556 29 1590
rect -29 1522 -17 1556
rect 17 1522 29 1556
rect -29 1483 29 1522
rect 129 2644 187 2683
rect 129 2610 141 2644
rect 175 2610 187 2644
rect 129 2576 187 2610
rect 129 2542 141 2576
rect 175 2542 187 2576
rect 129 2508 187 2542
rect 129 2474 141 2508
rect 175 2474 187 2508
rect 129 2440 187 2474
rect 129 2406 141 2440
rect 175 2406 187 2440
rect 129 2372 187 2406
rect 129 2338 141 2372
rect 175 2338 187 2372
rect 129 2304 187 2338
rect 129 2270 141 2304
rect 175 2270 187 2304
rect 129 2236 187 2270
rect 129 2202 141 2236
rect 175 2202 187 2236
rect 129 2168 187 2202
rect 129 2134 141 2168
rect 175 2134 187 2168
rect 129 2100 187 2134
rect 129 2066 141 2100
rect 175 2066 187 2100
rect 129 2032 187 2066
rect 129 1998 141 2032
rect 175 1998 187 2032
rect 129 1964 187 1998
rect 129 1930 141 1964
rect 175 1930 187 1964
rect 129 1896 187 1930
rect 129 1862 141 1896
rect 175 1862 187 1896
rect 129 1828 187 1862
rect 129 1794 141 1828
rect 175 1794 187 1828
rect 129 1760 187 1794
rect 129 1726 141 1760
rect 175 1726 187 1760
rect 129 1692 187 1726
rect 129 1658 141 1692
rect 175 1658 187 1692
rect 129 1624 187 1658
rect 129 1590 141 1624
rect 175 1590 187 1624
rect 129 1556 187 1590
rect 129 1522 141 1556
rect 175 1522 187 1556
rect 129 1483 187 1522
rect 287 2644 345 2683
rect 287 2610 299 2644
rect 333 2610 345 2644
rect 287 2576 345 2610
rect 287 2542 299 2576
rect 333 2542 345 2576
rect 287 2508 345 2542
rect 287 2474 299 2508
rect 333 2474 345 2508
rect 287 2440 345 2474
rect 287 2406 299 2440
rect 333 2406 345 2440
rect 287 2372 345 2406
rect 287 2338 299 2372
rect 333 2338 345 2372
rect 287 2304 345 2338
rect 287 2270 299 2304
rect 333 2270 345 2304
rect 287 2236 345 2270
rect 287 2202 299 2236
rect 333 2202 345 2236
rect 287 2168 345 2202
rect 287 2134 299 2168
rect 333 2134 345 2168
rect 287 2100 345 2134
rect 287 2066 299 2100
rect 333 2066 345 2100
rect 287 2032 345 2066
rect 287 1998 299 2032
rect 333 1998 345 2032
rect 287 1964 345 1998
rect 287 1930 299 1964
rect 333 1930 345 1964
rect 287 1896 345 1930
rect 287 1862 299 1896
rect 333 1862 345 1896
rect 287 1828 345 1862
rect 287 1794 299 1828
rect 333 1794 345 1828
rect 287 1760 345 1794
rect 287 1726 299 1760
rect 333 1726 345 1760
rect 287 1692 345 1726
rect 287 1658 299 1692
rect 333 1658 345 1692
rect 287 1624 345 1658
rect 287 1590 299 1624
rect 333 1590 345 1624
rect 287 1556 345 1590
rect 287 1522 299 1556
rect 333 1522 345 1556
rect 287 1483 345 1522
rect 445 2644 503 2683
rect 445 2610 457 2644
rect 491 2610 503 2644
rect 445 2576 503 2610
rect 445 2542 457 2576
rect 491 2542 503 2576
rect 445 2508 503 2542
rect 445 2474 457 2508
rect 491 2474 503 2508
rect 445 2440 503 2474
rect 445 2406 457 2440
rect 491 2406 503 2440
rect 445 2372 503 2406
rect 445 2338 457 2372
rect 491 2338 503 2372
rect 445 2304 503 2338
rect 445 2270 457 2304
rect 491 2270 503 2304
rect 445 2236 503 2270
rect 445 2202 457 2236
rect 491 2202 503 2236
rect 445 2168 503 2202
rect 445 2134 457 2168
rect 491 2134 503 2168
rect 445 2100 503 2134
rect 445 2066 457 2100
rect 491 2066 503 2100
rect 445 2032 503 2066
rect 445 1998 457 2032
rect 491 1998 503 2032
rect 445 1964 503 1998
rect 445 1930 457 1964
rect 491 1930 503 1964
rect 445 1896 503 1930
rect 445 1862 457 1896
rect 491 1862 503 1896
rect 445 1828 503 1862
rect 445 1794 457 1828
rect 491 1794 503 1828
rect 445 1760 503 1794
rect 445 1726 457 1760
rect 491 1726 503 1760
rect 445 1692 503 1726
rect 445 1658 457 1692
rect 491 1658 503 1692
rect 445 1624 503 1658
rect 445 1590 457 1624
rect 491 1590 503 1624
rect 445 1556 503 1590
rect 445 1522 457 1556
rect 491 1522 503 1556
rect 445 1483 503 1522
rect 603 2644 661 2683
rect 603 2610 615 2644
rect 649 2610 661 2644
rect 603 2576 661 2610
rect 603 2542 615 2576
rect 649 2542 661 2576
rect 603 2508 661 2542
rect 603 2474 615 2508
rect 649 2474 661 2508
rect 603 2440 661 2474
rect 603 2406 615 2440
rect 649 2406 661 2440
rect 603 2372 661 2406
rect 603 2338 615 2372
rect 649 2338 661 2372
rect 603 2304 661 2338
rect 603 2270 615 2304
rect 649 2270 661 2304
rect 603 2236 661 2270
rect 603 2202 615 2236
rect 649 2202 661 2236
rect 603 2168 661 2202
rect 603 2134 615 2168
rect 649 2134 661 2168
rect 603 2100 661 2134
rect 603 2066 615 2100
rect 649 2066 661 2100
rect 603 2032 661 2066
rect 603 1998 615 2032
rect 649 1998 661 2032
rect 603 1964 661 1998
rect 603 1930 615 1964
rect 649 1930 661 1964
rect 603 1896 661 1930
rect 603 1862 615 1896
rect 649 1862 661 1896
rect 603 1828 661 1862
rect 603 1794 615 1828
rect 649 1794 661 1828
rect 603 1760 661 1794
rect 603 1726 615 1760
rect 649 1726 661 1760
rect 603 1692 661 1726
rect 603 1658 615 1692
rect 649 1658 661 1692
rect 603 1624 661 1658
rect 603 1590 615 1624
rect 649 1590 661 1624
rect 603 1556 661 1590
rect 603 1522 615 1556
rect 649 1522 661 1556
rect 603 1483 661 1522
rect 761 2644 819 2683
rect 761 2610 773 2644
rect 807 2610 819 2644
rect 761 2576 819 2610
rect 761 2542 773 2576
rect 807 2542 819 2576
rect 761 2508 819 2542
rect 761 2474 773 2508
rect 807 2474 819 2508
rect 761 2440 819 2474
rect 761 2406 773 2440
rect 807 2406 819 2440
rect 761 2372 819 2406
rect 761 2338 773 2372
rect 807 2338 819 2372
rect 761 2304 819 2338
rect 761 2270 773 2304
rect 807 2270 819 2304
rect 761 2236 819 2270
rect 761 2202 773 2236
rect 807 2202 819 2236
rect 761 2168 819 2202
rect 761 2134 773 2168
rect 807 2134 819 2168
rect 761 2100 819 2134
rect 761 2066 773 2100
rect 807 2066 819 2100
rect 761 2032 819 2066
rect 761 1998 773 2032
rect 807 1998 819 2032
rect 761 1964 819 1998
rect 761 1930 773 1964
rect 807 1930 819 1964
rect 761 1896 819 1930
rect 761 1862 773 1896
rect 807 1862 819 1896
rect 761 1828 819 1862
rect 761 1794 773 1828
rect 807 1794 819 1828
rect 761 1760 819 1794
rect 761 1726 773 1760
rect 807 1726 819 1760
rect 761 1692 819 1726
rect 761 1658 773 1692
rect 807 1658 819 1692
rect 761 1624 819 1658
rect 761 1590 773 1624
rect 807 1590 819 1624
rect 761 1556 819 1590
rect 761 1522 773 1556
rect 807 1522 819 1556
rect 761 1483 819 1522
rect 919 2644 977 2683
rect 919 2610 931 2644
rect 965 2610 977 2644
rect 919 2576 977 2610
rect 919 2542 931 2576
rect 965 2542 977 2576
rect 919 2508 977 2542
rect 919 2474 931 2508
rect 965 2474 977 2508
rect 919 2440 977 2474
rect 919 2406 931 2440
rect 965 2406 977 2440
rect 919 2372 977 2406
rect 919 2338 931 2372
rect 965 2338 977 2372
rect 919 2304 977 2338
rect 919 2270 931 2304
rect 965 2270 977 2304
rect 919 2236 977 2270
rect 919 2202 931 2236
rect 965 2202 977 2236
rect 919 2168 977 2202
rect 919 2134 931 2168
rect 965 2134 977 2168
rect 919 2100 977 2134
rect 919 2066 931 2100
rect 965 2066 977 2100
rect 919 2032 977 2066
rect 919 1998 931 2032
rect 965 1998 977 2032
rect 919 1964 977 1998
rect 919 1930 931 1964
rect 965 1930 977 1964
rect 919 1896 977 1930
rect 919 1862 931 1896
rect 965 1862 977 1896
rect 919 1828 977 1862
rect 919 1794 931 1828
rect 965 1794 977 1828
rect 919 1760 977 1794
rect 919 1726 931 1760
rect 965 1726 977 1760
rect 919 1692 977 1726
rect 919 1658 931 1692
rect 965 1658 977 1692
rect 919 1624 977 1658
rect 919 1590 931 1624
rect 965 1590 977 1624
rect 919 1556 977 1590
rect 919 1522 931 1556
rect 965 1522 977 1556
rect 919 1483 977 1522
rect 1077 2644 1135 2683
rect 1077 2610 1089 2644
rect 1123 2610 1135 2644
rect 1077 2576 1135 2610
rect 1077 2542 1089 2576
rect 1123 2542 1135 2576
rect 1077 2508 1135 2542
rect 1077 2474 1089 2508
rect 1123 2474 1135 2508
rect 1077 2440 1135 2474
rect 1077 2406 1089 2440
rect 1123 2406 1135 2440
rect 1077 2372 1135 2406
rect 1077 2338 1089 2372
rect 1123 2338 1135 2372
rect 1077 2304 1135 2338
rect 1077 2270 1089 2304
rect 1123 2270 1135 2304
rect 1077 2236 1135 2270
rect 1077 2202 1089 2236
rect 1123 2202 1135 2236
rect 1077 2168 1135 2202
rect 1077 2134 1089 2168
rect 1123 2134 1135 2168
rect 1077 2100 1135 2134
rect 1077 2066 1089 2100
rect 1123 2066 1135 2100
rect 1077 2032 1135 2066
rect 1077 1998 1089 2032
rect 1123 1998 1135 2032
rect 1077 1964 1135 1998
rect 1077 1930 1089 1964
rect 1123 1930 1135 1964
rect 1077 1896 1135 1930
rect 1077 1862 1089 1896
rect 1123 1862 1135 1896
rect 1077 1828 1135 1862
rect 1077 1794 1089 1828
rect 1123 1794 1135 1828
rect 1077 1760 1135 1794
rect 1077 1726 1089 1760
rect 1123 1726 1135 1760
rect 1077 1692 1135 1726
rect 1077 1658 1089 1692
rect 1123 1658 1135 1692
rect 1077 1624 1135 1658
rect 1077 1590 1089 1624
rect 1123 1590 1135 1624
rect 1077 1556 1135 1590
rect 1077 1522 1089 1556
rect 1123 1522 1135 1556
rect 1077 1483 1135 1522
rect -1135 1279 -1077 1318
rect -1135 1245 -1123 1279
rect -1089 1245 -1077 1279
rect -1135 1211 -1077 1245
rect -1135 1177 -1123 1211
rect -1089 1177 -1077 1211
rect -1135 1143 -1077 1177
rect -1135 1109 -1123 1143
rect -1089 1109 -1077 1143
rect -1135 1075 -1077 1109
rect -1135 1041 -1123 1075
rect -1089 1041 -1077 1075
rect -1135 1007 -1077 1041
rect -1135 973 -1123 1007
rect -1089 973 -1077 1007
rect -1135 939 -1077 973
rect -1135 905 -1123 939
rect -1089 905 -1077 939
rect -1135 871 -1077 905
rect -1135 837 -1123 871
rect -1089 837 -1077 871
rect -1135 803 -1077 837
rect -1135 769 -1123 803
rect -1089 769 -1077 803
rect -1135 735 -1077 769
rect -1135 701 -1123 735
rect -1089 701 -1077 735
rect -1135 667 -1077 701
rect -1135 633 -1123 667
rect -1089 633 -1077 667
rect -1135 599 -1077 633
rect -1135 565 -1123 599
rect -1089 565 -1077 599
rect -1135 531 -1077 565
rect -1135 497 -1123 531
rect -1089 497 -1077 531
rect -1135 463 -1077 497
rect -1135 429 -1123 463
rect -1089 429 -1077 463
rect -1135 395 -1077 429
rect -1135 361 -1123 395
rect -1089 361 -1077 395
rect -1135 327 -1077 361
rect -1135 293 -1123 327
rect -1089 293 -1077 327
rect -1135 259 -1077 293
rect -1135 225 -1123 259
rect -1089 225 -1077 259
rect -1135 191 -1077 225
rect -1135 157 -1123 191
rect -1089 157 -1077 191
rect -1135 118 -1077 157
rect -977 1279 -919 1318
rect -977 1245 -965 1279
rect -931 1245 -919 1279
rect -977 1211 -919 1245
rect -977 1177 -965 1211
rect -931 1177 -919 1211
rect -977 1143 -919 1177
rect -977 1109 -965 1143
rect -931 1109 -919 1143
rect -977 1075 -919 1109
rect -977 1041 -965 1075
rect -931 1041 -919 1075
rect -977 1007 -919 1041
rect -977 973 -965 1007
rect -931 973 -919 1007
rect -977 939 -919 973
rect -977 905 -965 939
rect -931 905 -919 939
rect -977 871 -919 905
rect -977 837 -965 871
rect -931 837 -919 871
rect -977 803 -919 837
rect -977 769 -965 803
rect -931 769 -919 803
rect -977 735 -919 769
rect -977 701 -965 735
rect -931 701 -919 735
rect -977 667 -919 701
rect -977 633 -965 667
rect -931 633 -919 667
rect -977 599 -919 633
rect -977 565 -965 599
rect -931 565 -919 599
rect -977 531 -919 565
rect -977 497 -965 531
rect -931 497 -919 531
rect -977 463 -919 497
rect -977 429 -965 463
rect -931 429 -919 463
rect -977 395 -919 429
rect -977 361 -965 395
rect -931 361 -919 395
rect -977 327 -919 361
rect -977 293 -965 327
rect -931 293 -919 327
rect -977 259 -919 293
rect -977 225 -965 259
rect -931 225 -919 259
rect -977 191 -919 225
rect -977 157 -965 191
rect -931 157 -919 191
rect -977 118 -919 157
rect -819 1279 -761 1318
rect -819 1245 -807 1279
rect -773 1245 -761 1279
rect -819 1211 -761 1245
rect -819 1177 -807 1211
rect -773 1177 -761 1211
rect -819 1143 -761 1177
rect -819 1109 -807 1143
rect -773 1109 -761 1143
rect -819 1075 -761 1109
rect -819 1041 -807 1075
rect -773 1041 -761 1075
rect -819 1007 -761 1041
rect -819 973 -807 1007
rect -773 973 -761 1007
rect -819 939 -761 973
rect -819 905 -807 939
rect -773 905 -761 939
rect -819 871 -761 905
rect -819 837 -807 871
rect -773 837 -761 871
rect -819 803 -761 837
rect -819 769 -807 803
rect -773 769 -761 803
rect -819 735 -761 769
rect -819 701 -807 735
rect -773 701 -761 735
rect -819 667 -761 701
rect -819 633 -807 667
rect -773 633 -761 667
rect -819 599 -761 633
rect -819 565 -807 599
rect -773 565 -761 599
rect -819 531 -761 565
rect -819 497 -807 531
rect -773 497 -761 531
rect -819 463 -761 497
rect -819 429 -807 463
rect -773 429 -761 463
rect -819 395 -761 429
rect -819 361 -807 395
rect -773 361 -761 395
rect -819 327 -761 361
rect -819 293 -807 327
rect -773 293 -761 327
rect -819 259 -761 293
rect -819 225 -807 259
rect -773 225 -761 259
rect -819 191 -761 225
rect -819 157 -807 191
rect -773 157 -761 191
rect -819 118 -761 157
rect -661 1279 -603 1318
rect -661 1245 -649 1279
rect -615 1245 -603 1279
rect -661 1211 -603 1245
rect -661 1177 -649 1211
rect -615 1177 -603 1211
rect -661 1143 -603 1177
rect -661 1109 -649 1143
rect -615 1109 -603 1143
rect -661 1075 -603 1109
rect -661 1041 -649 1075
rect -615 1041 -603 1075
rect -661 1007 -603 1041
rect -661 973 -649 1007
rect -615 973 -603 1007
rect -661 939 -603 973
rect -661 905 -649 939
rect -615 905 -603 939
rect -661 871 -603 905
rect -661 837 -649 871
rect -615 837 -603 871
rect -661 803 -603 837
rect -661 769 -649 803
rect -615 769 -603 803
rect -661 735 -603 769
rect -661 701 -649 735
rect -615 701 -603 735
rect -661 667 -603 701
rect -661 633 -649 667
rect -615 633 -603 667
rect -661 599 -603 633
rect -661 565 -649 599
rect -615 565 -603 599
rect -661 531 -603 565
rect -661 497 -649 531
rect -615 497 -603 531
rect -661 463 -603 497
rect -661 429 -649 463
rect -615 429 -603 463
rect -661 395 -603 429
rect -661 361 -649 395
rect -615 361 -603 395
rect -661 327 -603 361
rect -661 293 -649 327
rect -615 293 -603 327
rect -661 259 -603 293
rect -661 225 -649 259
rect -615 225 -603 259
rect -661 191 -603 225
rect -661 157 -649 191
rect -615 157 -603 191
rect -661 118 -603 157
rect -503 1279 -445 1318
rect -503 1245 -491 1279
rect -457 1245 -445 1279
rect -503 1211 -445 1245
rect -503 1177 -491 1211
rect -457 1177 -445 1211
rect -503 1143 -445 1177
rect -503 1109 -491 1143
rect -457 1109 -445 1143
rect -503 1075 -445 1109
rect -503 1041 -491 1075
rect -457 1041 -445 1075
rect -503 1007 -445 1041
rect -503 973 -491 1007
rect -457 973 -445 1007
rect -503 939 -445 973
rect -503 905 -491 939
rect -457 905 -445 939
rect -503 871 -445 905
rect -503 837 -491 871
rect -457 837 -445 871
rect -503 803 -445 837
rect -503 769 -491 803
rect -457 769 -445 803
rect -503 735 -445 769
rect -503 701 -491 735
rect -457 701 -445 735
rect -503 667 -445 701
rect -503 633 -491 667
rect -457 633 -445 667
rect -503 599 -445 633
rect -503 565 -491 599
rect -457 565 -445 599
rect -503 531 -445 565
rect -503 497 -491 531
rect -457 497 -445 531
rect -503 463 -445 497
rect -503 429 -491 463
rect -457 429 -445 463
rect -503 395 -445 429
rect -503 361 -491 395
rect -457 361 -445 395
rect -503 327 -445 361
rect -503 293 -491 327
rect -457 293 -445 327
rect -503 259 -445 293
rect -503 225 -491 259
rect -457 225 -445 259
rect -503 191 -445 225
rect -503 157 -491 191
rect -457 157 -445 191
rect -503 118 -445 157
rect -345 1279 -287 1318
rect -345 1245 -333 1279
rect -299 1245 -287 1279
rect -345 1211 -287 1245
rect -345 1177 -333 1211
rect -299 1177 -287 1211
rect -345 1143 -287 1177
rect -345 1109 -333 1143
rect -299 1109 -287 1143
rect -345 1075 -287 1109
rect -345 1041 -333 1075
rect -299 1041 -287 1075
rect -345 1007 -287 1041
rect -345 973 -333 1007
rect -299 973 -287 1007
rect -345 939 -287 973
rect -345 905 -333 939
rect -299 905 -287 939
rect -345 871 -287 905
rect -345 837 -333 871
rect -299 837 -287 871
rect -345 803 -287 837
rect -345 769 -333 803
rect -299 769 -287 803
rect -345 735 -287 769
rect -345 701 -333 735
rect -299 701 -287 735
rect -345 667 -287 701
rect -345 633 -333 667
rect -299 633 -287 667
rect -345 599 -287 633
rect -345 565 -333 599
rect -299 565 -287 599
rect -345 531 -287 565
rect -345 497 -333 531
rect -299 497 -287 531
rect -345 463 -287 497
rect -345 429 -333 463
rect -299 429 -287 463
rect -345 395 -287 429
rect -345 361 -333 395
rect -299 361 -287 395
rect -345 327 -287 361
rect -345 293 -333 327
rect -299 293 -287 327
rect -345 259 -287 293
rect -345 225 -333 259
rect -299 225 -287 259
rect -345 191 -287 225
rect -345 157 -333 191
rect -299 157 -287 191
rect -345 118 -287 157
rect -187 1279 -129 1318
rect -187 1245 -175 1279
rect -141 1245 -129 1279
rect -187 1211 -129 1245
rect -187 1177 -175 1211
rect -141 1177 -129 1211
rect -187 1143 -129 1177
rect -187 1109 -175 1143
rect -141 1109 -129 1143
rect -187 1075 -129 1109
rect -187 1041 -175 1075
rect -141 1041 -129 1075
rect -187 1007 -129 1041
rect -187 973 -175 1007
rect -141 973 -129 1007
rect -187 939 -129 973
rect -187 905 -175 939
rect -141 905 -129 939
rect -187 871 -129 905
rect -187 837 -175 871
rect -141 837 -129 871
rect -187 803 -129 837
rect -187 769 -175 803
rect -141 769 -129 803
rect -187 735 -129 769
rect -187 701 -175 735
rect -141 701 -129 735
rect -187 667 -129 701
rect -187 633 -175 667
rect -141 633 -129 667
rect -187 599 -129 633
rect -187 565 -175 599
rect -141 565 -129 599
rect -187 531 -129 565
rect -187 497 -175 531
rect -141 497 -129 531
rect -187 463 -129 497
rect -187 429 -175 463
rect -141 429 -129 463
rect -187 395 -129 429
rect -187 361 -175 395
rect -141 361 -129 395
rect -187 327 -129 361
rect -187 293 -175 327
rect -141 293 -129 327
rect -187 259 -129 293
rect -187 225 -175 259
rect -141 225 -129 259
rect -187 191 -129 225
rect -187 157 -175 191
rect -141 157 -129 191
rect -187 118 -129 157
rect -29 1279 29 1318
rect -29 1245 -17 1279
rect 17 1245 29 1279
rect -29 1211 29 1245
rect -29 1177 -17 1211
rect 17 1177 29 1211
rect -29 1143 29 1177
rect -29 1109 -17 1143
rect 17 1109 29 1143
rect -29 1075 29 1109
rect -29 1041 -17 1075
rect 17 1041 29 1075
rect -29 1007 29 1041
rect -29 973 -17 1007
rect 17 973 29 1007
rect -29 939 29 973
rect -29 905 -17 939
rect 17 905 29 939
rect -29 871 29 905
rect -29 837 -17 871
rect 17 837 29 871
rect -29 803 29 837
rect -29 769 -17 803
rect 17 769 29 803
rect -29 735 29 769
rect -29 701 -17 735
rect 17 701 29 735
rect -29 667 29 701
rect -29 633 -17 667
rect 17 633 29 667
rect -29 599 29 633
rect -29 565 -17 599
rect 17 565 29 599
rect -29 531 29 565
rect -29 497 -17 531
rect 17 497 29 531
rect -29 463 29 497
rect -29 429 -17 463
rect 17 429 29 463
rect -29 395 29 429
rect -29 361 -17 395
rect 17 361 29 395
rect -29 327 29 361
rect -29 293 -17 327
rect 17 293 29 327
rect -29 259 29 293
rect -29 225 -17 259
rect 17 225 29 259
rect -29 191 29 225
rect -29 157 -17 191
rect 17 157 29 191
rect -29 118 29 157
rect 129 1279 187 1318
rect 129 1245 141 1279
rect 175 1245 187 1279
rect 129 1211 187 1245
rect 129 1177 141 1211
rect 175 1177 187 1211
rect 129 1143 187 1177
rect 129 1109 141 1143
rect 175 1109 187 1143
rect 129 1075 187 1109
rect 129 1041 141 1075
rect 175 1041 187 1075
rect 129 1007 187 1041
rect 129 973 141 1007
rect 175 973 187 1007
rect 129 939 187 973
rect 129 905 141 939
rect 175 905 187 939
rect 129 871 187 905
rect 129 837 141 871
rect 175 837 187 871
rect 129 803 187 837
rect 129 769 141 803
rect 175 769 187 803
rect 129 735 187 769
rect 129 701 141 735
rect 175 701 187 735
rect 129 667 187 701
rect 129 633 141 667
rect 175 633 187 667
rect 129 599 187 633
rect 129 565 141 599
rect 175 565 187 599
rect 129 531 187 565
rect 129 497 141 531
rect 175 497 187 531
rect 129 463 187 497
rect 129 429 141 463
rect 175 429 187 463
rect 129 395 187 429
rect 129 361 141 395
rect 175 361 187 395
rect 129 327 187 361
rect 129 293 141 327
rect 175 293 187 327
rect 129 259 187 293
rect 129 225 141 259
rect 175 225 187 259
rect 129 191 187 225
rect 129 157 141 191
rect 175 157 187 191
rect 129 118 187 157
rect 287 1279 345 1318
rect 287 1245 299 1279
rect 333 1245 345 1279
rect 287 1211 345 1245
rect 287 1177 299 1211
rect 333 1177 345 1211
rect 287 1143 345 1177
rect 287 1109 299 1143
rect 333 1109 345 1143
rect 287 1075 345 1109
rect 287 1041 299 1075
rect 333 1041 345 1075
rect 287 1007 345 1041
rect 287 973 299 1007
rect 333 973 345 1007
rect 287 939 345 973
rect 287 905 299 939
rect 333 905 345 939
rect 287 871 345 905
rect 287 837 299 871
rect 333 837 345 871
rect 287 803 345 837
rect 287 769 299 803
rect 333 769 345 803
rect 287 735 345 769
rect 287 701 299 735
rect 333 701 345 735
rect 287 667 345 701
rect 287 633 299 667
rect 333 633 345 667
rect 287 599 345 633
rect 287 565 299 599
rect 333 565 345 599
rect 287 531 345 565
rect 287 497 299 531
rect 333 497 345 531
rect 287 463 345 497
rect 287 429 299 463
rect 333 429 345 463
rect 287 395 345 429
rect 287 361 299 395
rect 333 361 345 395
rect 287 327 345 361
rect 287 293 299 327
rect 333 293 345 327
rect 287 259 345 293
rect 287 225 299 259
rect 333 225 345 259
rect 287 191 345 225
rect 287 157 299 191
rect 333 157 345 191
rect 287 118 345 157
rect 445 1279 503 1318
rect 445 1245 457 1279
rect 491 1245 503 1279
rect 445 1211 503 1245
rect 445 1177 457 1211
rect 491 1177 503 1211
rect 445 1143 503 1177
rect 445 1109 457 1143
rect 491 1109 503 1143
rect 445 1075 503 1109
rect 445 1041 457 1075
rect 491 1041 503 1075
rect 445 1007 503 1041
rect 445 973 457 1007
rect 491 973 503 1007
rect 445 939 503 973
rect 445 905 457 939
rect 491 905 503 939
rect 445 871 503 905
rect 445 837 457 871
rect 491 837 503 871
rect 445 803 503 837
rect 445 769 457 803
rect 491 769 503 803
rect 445 735 503 769
rect 445 701 457 735
rect 491 701 503 735
rect 445 667 503 701
rect 445 633 457 667
rect 491 633 503 667
rect 445 599 503 633
rect 445 565 457 599
rect 491 565 503 599
rect 445 531 503 565
rect 445 497 457 531
rect 491 497 503 531
rect 445 463 503 497
rect 445 429 457 463
rect 491 429 503 463
rect 445 395 503 429
rect 445 361 457 395
rect 491 361 503 395
rect 445 327 503 361
rect 445 293 457 327
rect 491 293 503 327
rect 445 259 503 293
rect 445 225 457 259
rect 491 225 503 259
rect 445 191 503 225
rect 445 157 457 191
rect 491 157 503 191
rect 445 118 503 157
rect 603 1279 661 1318
rect 603 1245 615 1279
rect 649 1245 661 1279
rect 603 1211 661 1245
rect 603 1177 615 1211
rect 649 1177 661 1211
rect 603 1143 661 1177
rect 603 1109 615 1143
rect 649 1109 661 1143
rect 603 1075 661 1109
rect 603 1041 615 1075
rect 649 1041 661 1075
rect 603 1007 661 1041
rect 603 973 615 1007
rect 649 973 661 1007
rect 603 939 661 973
rect 603 905 615 939
rect 649 905 661 939
rect 603 871 661 905
rect 603 837 615 871
rect 649 837 661 871
rect 603 803 661 837
rect 603 769 615 803
rect 649 769 661 803
rect 603 735 661 769
rect 603 701 615 735
rect 649 701 661 735
rect 603 667 661 701
rect 603 633 615 667
rect 649 633 661 667
rect 603 599 661 633
rect 603 565 615 599
rect 649 565 661 599
rect 603 531 661 565
rect 603 497 615 531
rect 649 497 661 531
rect 603 463 661 497
rect 603 429 615 463
rect 649 429 661 463
rect 603 395 661 429
rect 603 361 615 395
rect 649 361 661 395
rect 603 327 661 361
rect 603 293 615 327
rect 649 293 661 327
rect 603 259 661 293
rect 603 225 615 259
rect 649 225 661 259
rect 603 191 661 225
rect 603 157 615 191
rect 649 157 661 191
rect 603 118 661 157
rect 761 1279 819 1318
rect 761 1245 773 1279
rect 807 1245 819 1279
rect 761 1211 819 1245
rect 761 1177 773 1211
rect 807 1177 819 1211
rect 761 1143 819 1177
rect 761 1109 773 1143
rect 807 1109 819 1143
rect 761 1075 819 1109
rect 761 1041 773 1075
rect 807 1041 819 1075
rect 761 1007 819 1041
rect 761 973 773 1007
rect 807 973 819 1007
rect 761 939 819 973
rect 761 905 773 939
rect 807 905 819 939
rect 761 871 819 905
rect 761 837 773 871
rect 807 837 819 871
rect 761 803 819 837
rect 761 769 773 803
rect 807 769 819 803
rect 761 735 819 769
rect 761 701 773 735
rect 807 701 819 735
rect 761 667 819 701
rect 761 633 773 667
rect 807 633 819 667
rect 761 599 819 633
rect 761 565 773 599
rect 807 565 819 599
rect 761 531 819 565
rect 761 497 773 531
rect 807 497 819 531
rect 761 463 819 497
rect 761 429 773 463
rect 807 429 819 463
rect 761 395 819 429
rect 761 361 773 395
rect 807 361 819 395
rect 761 327 819 361
rect 761 293 773 327
rect 807 293 819 327
rect 761 259 819 293
rect 761 225 773 259
rect 807 225 819 259
rect 761 191 819 225
rect 761 157 773 191
rect 807 157 819 191
rect 761 118 819 157
rect 919 1279 977 1318
rect 919 1245 931 1279
rect 965 1245 977 1279
rect 919 1211 977 1245
rect 919 1177 931 1211
rect 965 1177 977 1211
rect 919 1143 977 1177
rect 919 1109 931 1143
rect 965 1109 977 1143
rect 919 1075 977 1109
rect 919 1041 931 1075
rect 965 1041 977 1075
rect 919 1007 977 1041
rect 919 973 931 1007
rect 965 973 977 1007
rect 919 939 977 973
rect 919 905 931 939
rect 965 905 977 939
rect 919 871 977 905
rect 919 837 931 871
rect 965 837 977 871
rect 919 803 977 837
rect 919 769 931 803
rect 965 769 977 803
rect 919 735 977 769
rect 919 701 931 735
rect 965 701 977 735
rect 919 667 977 701
rect 919 633 931 667
rect 965 633 977 667
rect 919 599 977 633
rect 919 565 931 599
rect 965 565 977 599
rect 919 531 977 565
rect 919 497 931 531
rect 965 497 977 531
rect 919 463 977 497
rect 919 429 931 463
rect 965 429 977 463
rect 919 395 977 429
rect 919 361 931 395
rect 965 361 977 395
rect 919 327 977 361
rect 919 293 931 327
rect 965 293 977 327
rect 919 259 977 293
rect 919 225 931 259
rect 965 225 977 259
rect 919 191 977 225
rect 919 157 931 191
rect 965 157 977 191
rect 919 118 977 157
rect 1077 1279 1135 1318
rect 1077 1245 1089 1279
rect 1123 1245 1135 1279
rect 1077 1211 1135 1245
rect 1077 1177 1089 1211
rect 1123 1177 1135 1211
rect 1077 1143 1135 1177
rect 1077 1109 1089 1143
rect 1123 1109 1135 1143
rect 1077 1075 1135 1109
rect 1077 1041 1089 1075
rect 1123 1041 1135 1075
rect 1077 1007 1135 1041
rect 1077 973 1089 1007
rect 1123 973 1135 1007
rect 1077 939 1135 973
rect 1077 905 1089 939
rect 1123 905 1135 939
rect 1077 871 1135 905
rect 1077 837 1089 871
rect 1123 837 1135 871
rect 1077 803 1135 837
rect 1077 769 1089 803
rect 1123 769 1135 803
rect 1077 735 1135 769
rect 1077 701 1089 735
rect 1123 701 1135 735
rect 1077 667 1135 701
rect 1077 633 1089 667
rect 1123 633 1135 667
rect 1077 599 1135 633
rect 1077 565 1089 599
rect 1123 565 1135 599
rect 1077 531 1135 565
rect 1077 497 1089 531
rect 1123 497 1135 531
rect 1077 463 1135 497
rect 1077 429 1089 463
rect 1123 429 1135 463
rect 1077 395 1135 429
rect 1077 361 1089 395
rect 1123 361 1135 395
rect 1077 327 1135 361
rect 1077 293 1089 327
rect 1123 293 1135 327
rect 1077 259 1135 293
rect 1077 225 1089 259
rect 1123 225 1135 259
rect 1077 191 1135 225
rect 1077 157 1089 191
rect 1123 157 1135 191
rect 1077 118 1135 157
rect -1135 -86 -1077 -47
rect -1135 -120 -1123 -86
rect -1089 -120 -1077 -86
rect -1135 -154 -1077 -120
rect -1135 -188 -1123 -154
rect -1089 -188 -1077 -154
rect -1135 -222 -1077 -188
rect -1135 -256 -1123 -222
rect -1089 -256 -1077 -222
rect -1135 -290 -1077 -256
rect -1135 -324 -1123 -290
rect -1089 -324 -1077 -290
rect -1135 -358 -1077 -324
rect -1135 -392 -1123 -358
rect -1089 -392 -1077 -358
rect -1135 -426 -1077 -392
rect -1135 -460 -1123 -426
rect -1089 -460 -1077 -426
rect -1135 -494 -1077 -460
rect -1135 -528 -1123 -494
rect -1089 -528 -1077 -494
rect -1135 -562 -1077 -528
rect -1135 -596 -1123 -562
rect -1089 -596 -1077 -562
rect -1135 -630 -1077 -596
rect -1135 -664 -1123 -630
rect -1089 -664 -1077 -630
rect -1135 -698 -1077 -664
rect -1135 -732 -1123 -698
rect -1089 -732 -1077 -698
rect -1135 -766 -1077 -732
rect -1135 -800 -1123 -766
rect -1089 -800 -1077 -766
rect -1135 -834 -1077 -800
rect -1135 -868 -1123 -834
rect -1089 -868 -1077 -834
rect -1135 -902 -1077 -868
rect -1135 -936 -1123 -902
rect -1089 -936 -1077 -902
rect -1135 -970 -1077 -936
rect -1135 -1004 -1123 -970
rect -1089 -1004 -1077 -970
rect -1135 -1038 -1077 -1004
rect -1135 -1072 -1123 -1038
rect -1089 -1072 -1077 -1038
rect -1135 -1106 -1077 -1072
rect -1135 -1140 -1123 -1106
rect -1089 -1140 -1077 -1106
rect -1135 -1174 -1077 -1140
rect -1135 -1208 -1123 -1174
rect -1089 -1208 -1077 -1174
rect -1135 -1247 -1077 -1208
rect -977 -86 -919 -47
rect -977 -120 -965 -86
rect -931 -120 -919 -86
rect -977 -154 -919 -120
rect -977 -188 -965 -154
rect -931 -188 -919 -154
rect -977 -222 -919 -188
rect -977 -256 -965 -222
rect -931 -256 -919 -222
rect -977 -290 -919 -256
rect -977 -324 -965 -290
rect -931 -324 -919 -290
rect -977 -358 -919 -324
rect -977 -392 -965 -358
rect -931 -392 -919 -358
rect -977 -426 -919 -392
rect -977 -460 -965 -426
rect -931 -460 -919 -426
rect -977 -494 -919 -460
rect -977 -528 -965 -494
rect -931 -528 -919 -494
rect -977 -562 -919 -528
rect -977 -596 -965 -562
rect -931 -596 -919 -562
rect -977 -630 -919 -596
rect -977 -664 -965 -630
rect -931 -664 -919 -630
rect -977 -698 -919 -664
rect -977 -732 -965 -698
rect -931 -732 -919 -698
rect -977 -766 -919 -732
rect -977 -800 -965 -766
rect -931 -800 -919 -766
rect -977 -834 -919 -800
rect -977 -868 -965 -834
rect -931 -868 -919 -834
rect -977 -902 -919 -868
rect -977 -936 -965 -902
rect -931 -936 -919 -902
rect -977 -970 -919 -936
rect -977 -1004 -965 -970
rect -931 -1004 -919 -970
rect -977 -1038 -919 -1004
rect -977 -1072 -965 -1038
rect -931 -1072 -919 -1038
rect -977 -1106 -919 -1072
rect -977 -1140 -965 -1106
rect -931 -1140 -919 -1106
rect -977 -1174 -919 -1140
rect -977 -1208 -965 -1174
rect -931 -1208 -919 -1174
rect -977 -1247 -919 -1208
rect -819 -86 -761 -47
rect -819 -120 -807 -86
rect -773 -120 -761 -86
rect -819 -154 -761 -120
rect -819 -188 -807 -154
rect -773 -188 -761 -154
rect -819 -222 -761 -188
rect -819 -256 -807 -222
rect -773 -256 -761 -222
rect -819 -290 -761 -256
rect -819 -324 -807 -290
rect -773 -324 -761 -290
rect -819 -358 -761 -324
rect -819 -392 -807 -358
rect -773 -392 -761 -358
rect -819 -426 -761 -392
rect -819 -460 -807 -426
rect -773 -460 -761 -426
rect -819 -494 -761 -460
rect -819 -528 -807 -494
rect -773 -528 -761 -494
rect -819 -562 -761 -528
rect -819 -596 -807 -562
rect -773 -596 -761 -562
rect -819 -630 -761 -596
rect -819 -664 -807 -630
rect -773 -664 -761 -630
rect -819 -698 -761 -664
rect -819 -732 -807 -698
rect -773 -732 -761 -698
rect -819 -766 -761 -732
rect -819 -800 -807 -766
rect -773 -800 -761 -766
rect -819 -834 -761 -800
rect -819 -868 -807 -834
rect -773 -868 -761 -834
rect -819 -902 -761 -868
rect -819 -936 -807 -902
rect -773 -936 -761 -902
rect -819 -970 -761 -936
rect -819 -1004 -807 -970
rect -773 -1004 -761 -970
rect -819 -1038 -761 -1004
rect -819 -1072 -807 -1038
rect -773 -1072 -761 -1038
rect -819 -1106 -761 -1072
rect -819 -1140 -807 -1106
rect -773 -1140 -761 -1106
rect -819 -1174 -761 -1140
rect -819 -1208 -807 -1174
rect -773 -1208 -761 -1174
rect -819 -1247 -761 -1208
rect -661 -86 -603 -47
rect -661 -120 -649 -86
rect -615 -120 -603 -86
rect -661 -154 -603 -120
rect -661 -188 -649 -154
rect -615 -188 -603 -154
rect -661 -222 -603 -188
rect -661 -256 -649 -222
rect -615 -256 -603 -222
rect -661 -290 -603 -256
rect -661 -324 -649 -290
rect -615 -324 -603 -290
rect -661 -358 -603 -324
rect -661 -392 -649 -358
rect -615 -392 -603 -358
rect -661 -426 -603 -392
rect -661 -460 -649 -426
rect -615 -460 -603 -426
rect -661 -494 -603 -460
rect -661 -528 -649 -494
rect -615 -528 -603 -494
rect -661 -562 -603 -528
rect -661 -596 -649 -562
rect -615 -596 -603 -562
rect -661 -630 -603 -596
rect -661 -664 -649 -630
rect -615 -664 -603 -630
rect -661 -698 -603 -664
rect -661 -732 -649 -698
rect -615 -732 -603 -698
rect -661 -766 -603 -732
rect -661 -800 -649 -766
rect -615 -800 -603 -766
rect -661 -834 -603 -800
rect -661 -868 -649 -834
rect -615 -868 -603 -834
rect -661 -902 -603 -868
rect -661 -936 -649 -902
rect -615 -936 -603 -902
rect -661 -970 -603 -936
rect -661 -1004 -649 -970
rect -615 -1004 -603 -970
rect -661 -1038 -603 -1004
rect -661 -1072 -649 -1038
rect -615 -1072 -603 -1038
rect -661 -1106 -603 -1072
rect -661 -1140 -649 -1106
rect -615 -1140 -603 -1106
rect -661 -1174 -603 -1140
rect -661 -1208 -649 -1174
rect -615 -1208 -603 -1174
rect -661 -1247 -603 -1208
rect -503 -86 -445 -47
rect -503 -120 -491 -86
rect -457 -120 -445 -86
rect -503 -154 -445 -120
rect -503 -188 -491 -154
rect -457 -188 -445 -154
rect -503 -222 -445 -188
rect -503 -256 -491 -222
rect -457 -256 -445 -222
rect -503 -290 -445 -256
rect -503 -324 -491 -290
rect -457 -324 -445 -290
rect -503 -358 -445 -324
rect -503 -392 -491 -358
rect -457 -392 -445 -358
rect -503 -426 -445 -392
rect -503 -460 -491 -426
rect -457 -460 -445 -426
rect -503 -494 -445 -460
rect -503 -528 -491 -494
rect -457 -528 -445 -494
rect -503 -562 -445 -528
rect -503 -596 -491 -562
rect -457 -596 -445 -562
rect -503 -630 -445 -596
rect -503 -664 -491 -630
rect -457 -664 -445 -630
rect -503 -698 -445 -664
rect -503 -732 -491 -698
rect -457 -732 -445 -698
rect -503 -766 -445 -732
rect -503 -800 -491 -766
rect -457 -800 -445 -766
rect -503 -834 -445 -800
rect -503 -868 -491 -834
rect -457 -868 -445 -834
rect -503 -902 -445 -868
rect -503 -936 -491 -902
rect -457 -936 -445 -902
rect -503 -970 -445 -936
rect -503 -1004 -491 -970
rect -457 -1004 -445 -970
rect -503 -1038 -445 -1004
rect -503 -1072 -491 -1038
rect -457 -1072 -445 -1038
rect -503 -1106 -445 -1072
rect -503 -1140 -491 -1106
rect -457 -1140 -445 -1106
rect -503 -1174 -445 -1140
rect -503 -1208 -491 -1174
rect -457 -1208 -445 -1174
rect -503 -1247 -445 -1208
rect -345 -86 -287 -47
rect -345 -120 -333 -86
rect -299 -120 -287 -86
rect -345 -154 -287 -120
rect -345 -188 -333 -154
rect -299 -188 -287 -154
rect -345 -222 -287 -188
rect -345 -256 -333 -222
rect -299 -256 -287 -222
rect -345 -290 -287 -256
rect -345 -324 -333 -290
rect -299 -324 -287 -290
rect -345 -358 -287 -324
rect -345 -392 -333 -358
rect -299 -392 -287 -358
rect -345 -426 -287 -392
rect -345 -460 -333 -426
rect -299 -460 -287 -426
rect -345 -494 -287 -460
rect -345 -528 -333 -494
rect -299 -528 -287 -494
rect -345 -562 -287 -528
rect -345 -596 -333 -562
rect -299 -596 -287 -562
rect -345 -630 -287 -596
rect -345 -664 -333 -630
rect -299 -664 -287 -630
rect -345 -698 -287 -664
rect -345 -732 -333 -698
rect -299 -732 -287 -698
rect -345 -766 -287 -732
rect -345 -800 -333 -766
rect -299 -800 -287 -766
rect -345 -834 -287 -800
rect -345 -868 -333 -834
rect -299 -868 -287 -834
rect -345 -902 -287 -868
rect -345 -936 -333 -902
rect -299 -936 -287 -902
rect -345 -970 -287 -936
rect -345 -1004 -333 -970
rect -299 -1004 -287 -970
rect -345 -1038 -287 -1004
rect -345 -1072 -333 -1038
rect -299 -1072 -287 -1038
rect -345 -1106 -287 -1072
rect -345 -1140 -333 -1106
rect -299 -1140 -287 -1106
rect -345 -1174 -287 -1140
rect -345 -1208 -333 -1174
rect -299 -1208 -287 -1174
rect -345 -1247 -287 -1208
rect -187 -86 -129 -47
rect -187 -120 -175 -86
rect -141 -120 -129 -86
rect -187 -154 -129 -120
rect -187 -188 -175 -154
rect -141 -188 -129 -154
rect -187 -222 -129 -188
rect -187 -256 -175 -222
rect -141 -256 -129 -222
rect -187 -290 -129 -256
rect -187 -324 -175 -290
rect -141 -324 -129 -290
rect -187 -358 -129 -324
rect -187 -392 -175 -358
rect -141 -392 -129 -358
rect -187 -426 -129 -392
rect -187 -460 -175 -426
rect -141 -460 -129 -426
rect -187 -494 -129 -460
rect -187 -528 -175 -494
rect -141 -528 -129 -494
rect -187 -562 -129 -528
rect -187 -596 -175 -562
rect -141 -596 -129 -562
rect -187 -630 -129 -596
rect -187 -664 -175 -630
rect -141 -664 -129 -630
rect -187 -698 -129 -664
rect -187 -732 -175 -698
rect -141 -732 -129 -698
rect -187 -766 -129 -732
rect -187 -800 -175 -766
rect -141 -800 -129 -766
rect -187 -834 -129 -800
rect -187 -868 -175 -834
rect -141 -868 -129 -834
rect -187 -902 -129 -868
rect -187 -936 -175 -902
rect -141 -936 -129 -902
rect -187 -970 -129 -936
rect -187 -1004 -175 -970
rect -141 -1004 -129 -970
rect -187 -1038 -129 -1004
rect -187 -1072 -175 -1038
rect -141 -1072 -129 -1038
rect -187 -1106 -129 -1072
rect -187 -1140 -175 -1106
rect -141 -1140 -129 -1106
rect -187 -1174 -129 -1140
rect -187 -1208 -175 -1174
rect -141 -1208 -129 -1174
rect -187 -1247 -129 -1208
rect -29 -86 29 -47
rect -29 -120 -17 -86
rect 17 -120 29 -86
rect -29 -154 29 -120
rect -29 -188 -17 -154
rect 17 -188 29 -154
rect -29 -222 29 -188
rect -29 -256 -17 -222
rect 17 -256 29 -222
rect -29 -290 29 -256
rect -29 -324 -17 -290
rect 17 -324 29 -290
rect -29 -358 29 -324
rect -29 -392 -17 -358
rect 17 -392 29 -358
rect -29 -426 29 -392
rect -29 -460 -17 -426
rect 17 -460 29 -426
rect -29 -494 29 -460
rect -29 -528 -17 -494
rect 17 -528 29 -494
rect -29 -562 29 -528
rect -29 -596 -17 -562
rect 17 -596 29 -562
rect -29 -630 29 -596
rect -29 -664 -17 -630
rect 17 -664 29 -630
rect -29 -698 29 -664
rect -29 -732 -17 -698
rect 17 -732 29 -698
rect -29 -766 29 -732
rect -29 -800 -17 -766
rect 17 -800 29 -766
rect -29 -834 29 -800
rect -29 -868 -17 -834
rect 17 -868 29 -834
rect -29 -902 29 -868
rect -29 -936 -17 -902
rect 17 -936 29 -902
rect -29 -970 29 -936
rect -29 -1004 -17 -970
rect 17 -1004 29 -970
rect -29 -1038 29 -1004
rect -29 -1072 -17 -1038
rect 17 -1072 29 -1038
rect -29 -1106 29 -1072
rect -29 -1140 -17 -1106
rect 17 -1140 29 -1106
rect -29 -1174 29 -1140
rect -29 -1208 -17 -1174
rect 17 -1208 29 -1174
rect -29 -1247 29 -1208
rect 129 -86 187 -47
rect 129 -120 141 -86
rect 175 -120 187 -86
rect 129 -154 187 -120
rect 129 -188 141 -154
rect 175 -188 187 -154
rect 129 -222 187 -188
rect 129 -256 141 -222
rect 175 -256 187 -222
rect 129 -290 187 -256
rect 129 -324 141 -290
rect 175 -324 187 -290
rect 129 -358 187 -324
rect 129 -392 141 -358
rect 175 -392 187 -358
rect 129 -426 187 -392
rect 129 -460 141 -426
rect 175 -460 187 -426
rect 129 -494 187 -460
rect 129 -528 141 -494
rect 175 -528 187 -494
rect 129 -562 187 -528
rect 129 -596 141 -562
rect 175 -596 187 -562
rect 129 -630 187 -596
rect 129 -664 141 -630
rect 175 -664 187 -630
rect 129 -698 187 -664
rect 129 -732 141 -698
rect 175 -732 187 -698
rect 129 -766 187 -732
rect 129 -800 141 -766
rect 175 -800 187 -766
rect 129 -834 187 -800
rect 129 -868 141 -834
rect 175 -868 187 -834
rect 129 -902 187 -868
rect 129 -936 141 -902
rect 175 -936 187 -902
rect 129 -970 187 -936
rect 129 -1004 141 -970
rect 175 -1004 187 -970
rect 129 -1038 187 -1004
rect 129 -1072 141 -1038
rect 175 -1072 187 -1038
rect 129 -1106 187 -1072
rect 129 -1140 141 -1106
rect 175 -1140 187 -1106
rect 129 -1174 187 -1140
rect 129 -1208 141 -1174
rect 175 -1208 187 -1174
rect 129 -1247 187 -1208
rect 287 -86 345 -47
rect 287 -120 299 -86
rect 333 -120 345 -86
rect 287 -154 345 -120
rect 287 -188 299 -154
rect 333 -188 345 -154
rect 287 -222 345 -188
rect 287 -256 299 -222
rect 333 -256 345 -222
rect 287 -290 345 -256
rect 287 -324 299 -290
rect 333 -324 345 -290
rect 287 -358 345 -324
rect 287 -392 299 -358
rect 333 -392 345 -358
rect 287 -426 345 -392
rect 287 -460 299 -426
rect 333 -460 345 -426
rect 287 -494 345 -460
rect 287 -528 299 -494
rect 333 -528 345 -494
rect 287 -562 345 -528
rect 287 -596 299 -562
rect 333 -596 345 -562
rect 287 -630 345 -596
rect 287 -664 299 -630
rect 333 -664 345 -630
rect 287 -698 345 -664
rect 287 -732 299 -698
rect 333 -732 345 -698
rect 287 -766 345 -732
rect 287 -800 299 -766
rect 333 -800 345 -766
rect 287 -834 345 -800
rect 287 -868 299 -834
rect 333 -868 345 -834
rect 287 -902 345 -868
rect 287 -936 299 -902
rect 333 -936 345 -902
rect 287 -970 345 -936
rect 287 -1004 299 -970
rect 333 -1004 345 -970
rect 287 -1038 345 -1004
rect 287 -1072 299 -1038
rect 333 -1072 345 -1038
rect 287 -1106 345 -1072
rect 287 -1140 299 -1106
rect 333 -1140 345 -1106
rect 287 -1174 345 -1140
rect 287 -1208 299 -1174
rect 333 -1208 345 -1174
rect 287 -1247 345 -1208
rect 445 -86 503 -47
rect 445 -120 457 -86
rect 491 -120 503 -86
rect 445 -154 503 -120
rect 445 -188 457 -154
rect 491 -188 503 -154
rect 445 -222 503 -188
rect 445 -256 457 -222
rect 491 -256 503 -222
rect 445 -290 503 -256
rect 445 -324 457 -290
rect 491 -324 503 -290
rect 445 -358 503 -324
rect 445 -392 457 -358
rect 491 -392 503 -358
rect 445 -426 503 -392
rect 445 -460 457 -426
rect 491 -460 503 -426
rect 445 -494 503 -460
rect 445 -528 457 -494
rect 491 -528 503 -494
rect 445 -562 503 -528
rect 445 -596 457 -562
rect 491 -596 503 -562
rect 445 -630 503 -596
rect 445 -664 457 -630
rect 491 -664 503 -630
rect 445 -698 503 -664
rect 445 -732 457 -698
rect 491 -732 503 -698
rect 445 -766 503 -732
rect 445 -800 457 -766
rect 491 -800 503 -766
rect 445 -834 503 -800
rect 445 -868 457 -834
rect 491 -868 503 -834
rect 445 -902 503 -868
rect 445 -936 457 -902
rect 491 -936 503 -902
rect 445 -970 503 -936
rect 445 -1004 457 -970
rect 491 -1004 503 -970
rect 445 -1038 503 -1004
rect 445 -1072 457 -1038
rect 491 -1072 503 -1038
rect 445 -1106 503 -1072
rect 445 -1140 457 -1106
rect 491 -1140 503 -1106
rect 445 -1174 503 -1140
rect 445 -1208 457 -1174
rect 491 -1208 503 -1174
rect 445 -1247 503 -1208
rect 603 -86 661 -47
rect 603 -120 615 -86
rect 649 -120 661 -86
rect 603 -154 661 -120
rect 603 -188 615 -154
rect 649 -188 661 -154
rect 603 -222 661 -188
rect 603 -256 615 -222
rect 649 -256 661 -222
rect 603 -290 661 -256
rect 603 -324 615 -290
rect 649 -324 661 -290
rect 603 -358 661 -324
rect 603 -392 615 -358
rect 649 -392 661 -358
rect 603 -426 661 -392
rect 603 -460 615 -426
rect 649 -460 661 -426
rect 603 -494 661 -460
rect 603 -528 615 -494
rect 649 -528 661 -494
rect 603 -562 661 -528
rect 603 -596 615 -562
rect 649 -596 661 -562
rect 603 -630 661 -596
rect 603 -664 615 -630
rect 649 -664 661 -630
rect 603 -698 661 -664
rect 603 -732 615 -698
rect 649 -732 661 -698
rect 603 -766 661 -732
rect 603 -800 615 -766
rect 649 -800 661 -766
rect 603 -834 661 -800
rect 603 -868 615 -834
rect 649 -868 661 -834
rect 603 -902 661 -868
rect 603 -936 615 -902
rect 649 -936 661 -902
rect 603 -970 661 -936
rect 603 -1004 615 -970
rect 649 -1004 661 -970
rect 603 -1038 661 -1004
rect 603 -1072 615 -1038
rect 649 -1072 661 -1038
rect 603 -1106 661 -1072
rect 603 -1140 615 -1106
rect 649 -1140 661 -1106
rect 603 -1174 661 -1140
rect 603 -1208 615 -1174
rect 649 -1208 661 -1174
rect 603 -1247 661 -1208
rect 761 -86 819 -47
rect 761 -120 773 -86
rect 807 -120 819 -86
rect 761 -154 819 -120
rect 761 -188 773 -154
rect 807 -188 819 -154
rect 761 -222 819 -188
rect 761 -256 773 -222
rect 807 -256 819 -222
rect 761 -290 819 -256
rect 761 -324 773 -290
rect 807 -324 819 -290
rect 761 -358 819 -324
rect 761 -392 773 -358
rect 807 -392 819 -358
rect 761 -426 819 -392
rect 761 -460 773 -426
rect 807 -460 819 -426
rect 761 -494 819 -460
rect 761 -528 773 -494
rect 807 -528 819 -494
rect 761 -562 819 -528
rect 761 -596 773 -562
rect 807 -596 819 -562
rect 761 -630 819 -596
rect 761 -664 773 -630
rect 807 -664 819 -630
rect 761 -698 819 -664
rect 761 -732 773 -698
rect 807 -732 819 -698
rect 761 -766 819 -732
rect 761 -800 773 -766
rect 807 -800 819 -766
rect 761 -834 819 -800
rect 761 -868 773 -834
rect 807 -868 819 -834
rect 761 -902 819 -868
rect 761 -936 773 -902
rect 807 -936 819 -902
rect 761 -970 819 -936
rect 761 -1004 773 -970
rect 807 -1004 819 -970
rect 761 -1038 819 -1004
rect 761 -1072 773 -1038
rect 807 -1072 819 -1038
rect 761 -1106 819 -1072
rect 761 -1140 773 -1106
rect 807 -1140 819 -1106
rect 761 -1174 819 -1140
rect 761 -1208 773 -1174
rect 807 -1208 819 -1174
rect 761 -1247 819 -1208
rect 919 -86 977 -47
rect 919 -120 931 -86
rect 965 -120 977 -86
rect 919 -154 977 -120
rect 919 -188 931 -154
rect 965 -188 977 -154
rect 919 -222 977 -188
rect 919 -256 931 -222
rect 965 -256 977 -222
rect 919 -290 977 -256
rect 919 -324 931 -290
rect 965 -324 977 -290
rect 919 -358 977 -324
rect 919 -392 931 -358
rect 965 -392 977 -358
rect 919 -426 977 -392
rect 919 -460 931 -426
rect 965 -460 977 -426
rect 919 -494 977 -460
rect 919 -528 931 -494
rect 965 -528 977 -494
rect 919 -562 977 -528
rect 919 -596 931 -562
rect 965 -596 977 -562
rect 919 -630 977 -596
rect 919 -664 931 -630
rect 965 -664 977 -630
rect 919 -698 977 -664
rect 919 -732 931 -698
rect 965 -732 977 -698
rect 919 -766 977 -732
rect 919 -800 931 -766
rect 965 -800 977 -766
rect 919 -834 977 -800
rect 919 -868 931 -834
rect 965 -868 977 -834
rect 919 -902 977 -868
rect 919 -936 931 -902
rect 965 -936 977 -902
rect 919 -970 977 -936
rect 919 -1004 931 -970
rect 965 -1004 977 -970
rect 919 -1038 977 -1004
rect 919 -1072 931 -1038
rect 965 -1072 977 -1038
rect 919 -1106 977 -1072
rect 919 -1140 931 -1106
rect 965 -1140 977 -1106
rect 919 -1174 977 -1140
rect 919 -1208 931 -1174
rect 965 -1208 977 -1174
rect 919 -1247 977 -1208
rect 1077 -86 1135 -47
rect 1077 -120 1089 -86
rect 1123 -120 1135 -86
rect 1077 -154 1135 -120
rect 1077 -188 1089 -154
rect 1123 -188 1135 -154
rect 1077 -222 1135 -188
rect 1077 -256 1089 -222
rect 1123 -256 1135 -222
rect 1077 -290 1135 -256
rect 1077 -324 1089 -290
rect 1123 -324 1135 -290
rect 1077 -358 1135 -324
rect 1077 -392 1089 -358
rect 1123 -392 1135 -358
rect 1077 -426 1135 -392
rect 1077 -460 1089 -426
rect 1123 -460 1135 -426
rect 1077 -494 1135 -460
rect 1077 -528 1089 -494
rect 1123 -528 1135 -494
rect 1077 -562 1135 -528
rect 1077 -596 1089 -562
rect 1123 -596 1135 -562
rect 1077 -630 1135 -596
rect 1077 -664 1089 -630
rect 1123 -664 1135 -630
rect 1077 -698 1135 -664
rect 1077 -732 1089 -698
rect 1123 -732 1135 -698
rect 1077 -766 1135 -732
rect 1077 -800 1089 -766
rect 1123 -800 1135 -766
rect 1077 -834 1135 -800
rect 1077 -868 1089 -834
rect 1123 -868 1135 -834
rect 1077 -902 1135 -868
rect 1077 -936 1089 -902
rect 1123 -936 1135 -902
rect 1077 -970 1135 -936
rect 1077 -1004 1089 -970
rect 1123 -1004 1135 -970
rect 1077 -1038 1135 -1004
rect 1077 -1072 1089 -1038
rect 1123 -1072 1135 -1038
rect 1077 -1106 1135 -1072
rect 1077 -1140 1089 -1106
rect 1123 -1140 1135 -1106
rect 1077 -1174 1135 -1140
rect 1077 -1208 1089 -1174
rect 1123 -1208 1135 -1174
rect 1077 -1247 1135 -1208
rect -1135 -1451 -1077 -1412
rect -1135 -1485 -1123 -1451
rect -1089 -1485 -1077 -1451
rect -1135 -1519 -1077 -1485
rect -1135 -1553 -1123 -1519
rect -1089 -1553 -1077 -1519
rect -1135 -1587 -1077 -1553
rect -1135 -1621 -1123 -1587
rect -1089 -1621 -1077 -1587
rect -1135 -1655 -1077 -1621
rect -1135 -1689 -1123 -1655
rect -1089 -1689 -1077 -1655
rect -1135 -1723 -1077 -1689
rect -1135 -1757 -1123 -1723
rect -1089 -1757 -1077 -1723
rect -1135 -1791 -1077 -1757
rect -1135 -1825 -1123 -1791
rect -1089 -1825 -1077 -1791
rect -1135 -1859 -1077 -1825
rect -1135 -1893 -1123 -1859
rect -1089 -1893 -1077 -1859
rect -1135 -1927 -1077 -1893
rect -1135 -1961 -1123 -1927
rect -1089 -1961 -1077 -1927
rect -1135 -1995 -1077 -1961
rect -1135 -2029 -1123 -1995
rect -1089 -2029 -1077 -1995
rect -1135 -2063 -1077 -2029
rect -1135 -2097 -1123 -2063
rect -1089 -2097 -1077 -2063
rect -1135 -2131 -1077 -2097
rect -1135 -2165 -1123 -2131
rect -1089 -2165 -1077 -2131
rect -1135 -2199 -1077 -2165
rect -1135 -2233 -1123 -2199
rect -1089 -2233 -1077 -2199
rect -1135 -2267 -1077 -2233
rect -1135 -2301 -1123 -2267
rect -1089 -2301 -1077 -2267
rect -1135 -2335 -1077 -2301
rect -1135 -2369 -1123 -2335
rect -1089 -2369 -1077 -2335
rect -1135 -2403 -1077 -2369
rect -1135 -2437 -1123 -2403
rect -1089 -2437 -1077 -2403
rect -1135 -2471 -1077 -2437
rect -1135 -2505 -1123 -2471
rect -1089 -2505 -1077 -2471
rect -1135 -2539 -1077 -2505
rect -1135 -2573 -1123 -2539
rect -1089 -2573 -1077 -2539
rect -1135 -2612 -1077 -2573
rect -977 -1451 -919 -1412
rect -977 -1485 -965 -1451
rect -931 -1485 -919 -1451
rect -977 -1519 -919 -1485
rect -977 -1553 -965 -1519
rect -931 -1553 -919 -1519
rect -977 -1587 -919 -1553
rect -977 -1621 -965 -1587
rect -931 -1621 -919 -1587
rect -977 -1655 -919 -1621
rect -977 -1689 -965 -1655
rect -931 -1689 -919 -1655
rect -977 -1723 -919 -1689
rect -977 -1757 -965 -1723
rect -931 -1757 -919 -1723
rect -977 -1791 -919 -1757
rect -977 -1825 -965 -1791
rect -931 -1825 -919 -1791
rect -977 -1859 -919 -1825
rect -977 -1893 -965 -1859
rect -931 -1893 -919 -1859
rect -977 -1927 -919 -1893
rect -977 -1961 -965 -1927
rect -931 -1961 -919 -1927
rect -977 -1995 -919 -1961
rect -977 -2029 -965 -1995
rect -931 -2029 -919 -1995
rect -977 -2063 -919 -2029
rect -977 -2097 -965 -2063
rect -931 -2097 -919 -2063
rect -977 -2131 -919 -2097
rect -977 -2165 -965 -2131
rect -931 -2165 -919 -2131
rect -977 -2199 -919 -2165
rect -977 -2233 -965 -2199
rect -931 -2233 -919 -2199
rect -977 -2267 -919 -2233
rect -977 -2301 -965 -2267
rect -931 -2301 -919 -2267
rect -977 -2335 -919 -2301
rect -977 -2369 -965 -2335
rect -931 -2369 -919 -2335
rect -977 -2403 -919 -2369
rect -977 -2437 -965 -2403
rect -931 -2437 -919 -2403
rect -977 -2471 -919 -2437
rect -977 -2505 -965 -2471
rect -931 -2505 -919 -2471
rect -977 -2539 -919 -2505
rect -977 -2573 -965 -2539
rect -931 -2573 -919 -2539
rect -977 -2612 -919 -2573
rect -819 -1451 -761 -1412
rect -819 -1485 -807 -1451
rect -773 -1485 -761 -1451
rect -819 -1519 -761 -1485
rect -819 -1553 -807 -1519
rect -773 -1553 -761 -1519
rect -819 -1587 -761 -1553
rect -819 -1621 -807 -1587
rect -773 -1621 -761 -1587
rect -819 -1655 -761 -1621
rect -819 -1689 -807 -1655
rect -773 -1689 -761 -1655
rect -819 -1723 -761 -1689
rect -819 -1757 -807 -1723
rect -773 -1757 -761 -1723
rect -819 -1791 -761 -1757
rect -819 -1825 -807 -1791
rect -773 -1825 -761 -1791
rect -819 -1859 -761 -1825
rect -819 -1893 -807 -1859
rect -773 -1893 -761 -1859
rect -819 -1927 -761 -1893
rect -819 -1961 -807 -1927
rect -773 -1961 -761 -1927
rect -819 -1995 -761 -1961
rect -819 -2029 -807 -1995
rect -773 -2029 -761 -1995
rect -819 -2063 -761 -2029
rect -819 -2097 -807 -2063
rect -773 -2097 -761 -2063
rect -819 -2131 -761 -2097
rect -819 -2165 -807 -2131
rect -773 -2165 -761 -2131
rect -819 -2199 -761 -2165
rect -819 -2233 -807 -2199
rect -773 -2233 -761 -2199
rect -819 -2267 -761 -2233
rect -819 -2301 -807 -2267
rect -773 -2301 -761 -2267
rect -819 -2335 -761 -2301
rect -819 -2369 -807 -2335
rect -773 -2369 -761 -2335
rect -819 -2403 -761 -2369
rect -819 -2437 -807 -2403
rect -773 -2437 -761 -2403
rect -819 -2471 -761 -2437
rect -819 -2505 -807 -2471
rect -773 -2505 -761 -2471
rect -819 -2539 -761 -2505
rect -819 -2573 -807 -2539
rect -773 -2573 -761 -2539
rect -819 -2612 -761 -2573
rect -661 -1451 -603 -1412
rect -661 -1485 -649 -1451
rect -615 -1485 -603 -1451
rect -661 -1519 -603 -1485
rect -661 -1553 -649 -1519
rect -615 -1553 -603 -1519
rect -661 -1587 -603 -1553
rect -661 -1621 -649 -1587
rect -615 -1621 -603 -1587
rect -661 -1655 -603 -1621
rect -661 -1689 -649 -1655
rect -615 -1689 -603 -1655
rect -661 -1723 -603 -1689
rect -661 -1757 -649 -1723
rect -615 -1757 -603 -1723
rect -661 -1791 -603 -1757
rect -661 -1825 -649 -1791
rect -615 -1825 -603 -1791
rect -661 -1859 -603 -1825
rect -661 -1893 -649 -1859
rect -615 -1893 -603 -1859
rect -661 -1927 -603 -1893
rect -661 -1961 -649 -1927
rect -615 -1961 -603 -1927
rect -661 -1995 -603 -1961
rect -661 -2029 -649 -1995
rect -615 -2029 -603 -1995
rect -661 -2063 -603 -2029
rect -661 -2097 -649 -2063
rect -615 -2097 -603 -2063
rect -661 -2131 -603 -2097
rect -661 -2165 -649 -2131
rect -615 -2165 -603 -2131
rect -661 -2199 -603 -2165
rect -661 -2233 -649 -2199
rect -615 -2233 -603 -2199
rect -661 -2267 -603 -2233
rect -661 -2301 -649 -2267
rect -615 -2301 -603 -2267
rect -661 -2335 -603 -2301
rect -661 -2369 -649 -2335
rect -615 -2369 -603 -2335
rect -661 -2403 -603 -2369
rect -661 -2437 -649 -2403
rect -615 -2437 -603 -2403
rect -661 -2471 -603 -2437
rect -661 -2505 -649 -2471
rect -615 -2505 -603 -2471
rect -661 -2539 -603 -2505
rect -661 -2573 -649 -2539
rect -615 -2573 -603 -2539
rect -661 -2612 -603 -2573
rect -503 -1451 -445 -1412
rect -503 -1485 -491 -1451
rect -457 -1485 -445 -1451
rect -503 -1519 -445 -1485
rect -503 -1553 -491 -1519
rect -457 -1553 -445 -1519
rect -503 -1587 -445 -1553
rect -503 -1621 -491 -1587
rect -457 -1621 -445 -1587
rect -503 -1655 -445 -1621
rect -503 -1689 -491 -1655
rect -457 -1689 -445 -1655
rect -503 -1723 -445 -1689
rect -503 -1757 -491 -1723
rect -457 -1757 -445 -1723
rect -503 -1791 -445 -1757
rect -503 -1825 -491 -1791
rect -457 -1825 -445 -1791
rect -503 -1859 -445 -1825
rect -503 -1893 -491 -1859
rect -457 -1893 -445 -1859
rect -503 -1927 -445 -1893
rect -503 -1961 -491 -1927
rect -457 -1961 -445 -1927
rect -503 -1995 -445 -1961
rect -503 -2029 -491 -1995
rect -457 -2029 -445 -1995
rect -503 -2063 -445 -2029
rect -503 -2097 -491 -2063
rect -457 -2097 -445 -2063
rect -503 -2131 -445 -2097
rect -503 -2165 -491 -2131
rect -457 -2165 -445 -2131
rect -503 -2199 -445 -2165
rect -503 -2233 -491 -2199
rect -457 -2233 -445 -2199
rect -503 -2267 -445 -2233
rect -503 -2301 -491 -2267
rect -457 -2301 -445 -2267
rect -503 -2335 -445 -2301
rect -503 -2369 -491 -2335
rect -457 -2369 -445 -2335
rect -503 -2403 -445 -2369
rect -503 -2437 -491 -2403
rect -457 -2437 -445 -2403
rect -503 -2471 -445 -2437
rect -503 -2505 -491 -2471
rect -457 -2505 -445 -2471
rect -503 -2539 -445 -2505
rect -503 -2573 -491 -2539
rect -457 -2573 -445 -2539
rect -503 -2612 -445 -2573
rect -345 -1451 -287 -1412
rect -345 -1485 -333 -1451
rect -299 -1485 -287 -1451
rect -345 -1519 -287 -1485
rect -345 -1553 -333 -1519
rect -299 -1553 -287 -1519
rect -345 -1587 -287 -1553
rect -345 -1621 -333 -1587
rect -299 -1621 -287 -1587
rect -345 -1655 -287 -1621
rect -345 -1689 -333 -1655
rect -299 -1689 -287 -1655
rect -345 -1723 -287 -1689
rect -345 -1757 -333 -1723
rect -299 -1757 -287 -1723
rect -345 -1791 -287 -1757
rect -345 -1825 -333 -1791
rect -299 -1825 -287 -1791
rect -345 -1859 -287 -1825
rect -345 -1893 -333 -1859
rect -299 -1893 -287 -1859
rect -345 -1927 -287 -1893
rect -345 -1961 -333 -1927
rect -299 -1961 -287 -1927
rect -345 -1995 -287 -1961
rect -345 -2029 -333 -1995
rect -299 -2029 -287 -1995
rect -345 -2063 -287 -2029
rect -345 -2097 -333 -2063
rect -299 -2097 -287 -2063
rect -345 -2131 -287 -2097
rect -345 -2165 -333 -2131
rect -299 -2165 -287 -2131
rect -345 -2199 -287 -2165
rect -345 -2233 -333 -2199
rect -299 -2233 -287 -2199
rect -345 -2267 -287 -2233
rect -345 -2301 -333 -2267
rect -299 -2301 -287 -2267
rect -345 -2335 -287 -2301
rect -345 -2369 -333 -2335
rect -299 -2369 -287 -2335
rect -345 -2403 -287 -2369
rect -345 -2437 -333 -2403
rect -299 -2437 -287 -2403
rect -345 -2471 -287 -2437
rect -345 -2505 -333 -2471
rect -299 -2505 -287 -2471
rect -345 -2539 -287 -2505
rect -345 -2573 -333 -2539
rect -299 -2573 -287 -2539
rect -345 -2612 -287 -2573
rect -187 -1451 -129 -1412
rect -187 -1485 -175 -1451
rect -141 -1485 -129 -1451
rect -187 -1519 -129 -1485
rect -187 -1553 -175 -1519
rect -141 -1553 -129 -1519
rect -187 -1587 -129 -1553
rect -187 -1621 -175 -1587
rect -141 -1621 -129 -1587
rect -187 -1655 -129 -1621
rect -187 -1689 -175 -1655
rect -141 -1689 -129 -1655
rect -187 -1723 -129 -1689
rect -187 -1757 -175 -1723
rect -141 -1757 -129 -1723
rect -187 -1791 -129 -1757
rect -187 -1825 -175 -1791
rect -141 -1825 -129 -1791
rect -187 -1859 -129 -1825
rect -187 -1893 -175 -1859
rect -141 -1893 -129 -1859
rect -187 -1927 -129 -1893
rect -187 -1961 -175 -1927
rect -141 -1961 -129 -1927
rect -187 -1995 -129 -1961
rect -187 -2029 -175 -1995
rect -141 -2029 -129 -1995
rect -187 -2063 -129 -2029
rect -187 -2097 -175 -2063
rect -141 -2097 -129 -2063
rect -187 -2131 -129 -2097
rect -187 -2165 -175 -2131
rect -141 -2165 -129 -2131
rect -187 -2199 -129 -2165
rect -187 -2233 -175 -2199
rect -141 -2233 -129 -2199
rect -187 -2267 -129 -2233
rect -187 -2301 -175 -2267
rect -141 -2301 -129 -2267
rect -187 -2335 -129 -2301
rect -187 -2369 -175 -2335
rect -141 -2369 -129 -2335
rect -187 -2403 -129 -2369
rect -187 -2437 -175 -2403
rect -141 -2437 -129 -2403
rect -187 -2471 -129 -2437
rect -187 -2505 -175 -2471
rect -141 -2505 -129 -2471
rect -187 -2539 -129 -2505
rect -187 -2573 -175 -2539
rect -141 -2573 -129 -2539
rect -187 -2612 -129 -2573
rect -29 -1451 29 -1412
rect -29 -1485 -17 -1451
rect 17 -1485 29 -1451
rect -29 -1519 29 -1485
rect -29 -1553 -17 -1519
rect 17 -1553 29 -1519
rect -29 -1587 29 -1553
rect -29 -1621 -17 -1587
rect 17 -1621 29 -1587
rect -29 -1655 29 -1621
rect -29 -1689 -17 -1655
rect 17 -1689 29 -1655
rect -29 -1723 29 -1689
rect -29 -1757 -17 -1723
rect 17 -1757 29 -1723
rect -29 -1791 29 -1757
rect -29 -1825 -17 -1791
rect 17 -1825 29 -1791
rect -29 -1859 29 -1825
rect -29 -1893 -17 -1859
rect 17 -1893 29 -1859
rect -29 -1927 29 -1893
rect -29 -1961 -17 -1927
rect 17 -1961 29 -1927
rect -29 -1995 29 -1961
rect -29 -2029 -17 -1995
rect 17 -2029 29 -1995
rect -29 -2063 29 -2029
rect -29 -2097 -17 -2063
rect 17 -2097 29 -2063
rect -29 -2131 29 -2097
rect -29 -2165 -17 -2131
rect 17 -2165 29 -2131
rect -29 -2199 29 -2165
rect -29 -2233 -17 -2199
rect 17 -2233 29 -2199
rect -29 -2267 29 -2233
rect -29 -2301 -17 -2267
rect 17 -2301 29 -2267
rect -29 -2335 29 -2301
rect -29 -2369 -17 -2335
rect 17 -2369 29 -2335
rect -29 -2403 29 -2369
rect -29 -2437 -17 -2403
rect 17 -2437 29 -2403
rect -29 -2471 29 -2437
rect -29 -2505 -17 -2471
rect 17 -2505 29 -2471
rect -29 -2539 29 -2505
rect -29 -2573 -17 -2539
rect 17 -2573 29 -2539
rect -29 -2612 29 -2573
rect 129 -1451 187 -1412
rect 129 -1485 141 -1451
rect 175 -1485 187 -1451
rect 129 -1519 187 -1485
rect 129 -1553 141 -1519
rect 175 -1553 187 -1519
rect 129 -1587 187 -1553
rect 129 -1621 141 -1587
rect 175 -1621 187 -1587
rect 129 -1655 187 -1621
rect 129 -1689 141 -1655
rect 175 -1689 187 -1655
rect 129 -1723 187 -1689
rect 129 -1757 141 -1723
rect 175 -1757 187 -1723
rect 129 -1791 187 -1757
rect 129 -1825 141 -1791
rect 175 -1825 187 -1791
rect 129 -1859 187 -1825
rect 129 -1893 141 -1859
rect 175 -1893 187 -1859
rect 129 -1927 187 -1893
rect 129 -1961 141 -1927
rect 175 -1961 187 -1927
rect 129 -1995 187 -1961
rect 129 -2029 141 -1995
rect 175 -2029 187 -1995
rect 129 -2063 187 -2029
rect 129 -2097 141 -2063
rect 175 -2097 187 -2063
rect 129 -2131 187 -2097
rect 129 -2165 141 -2131
rect 175 -2165 187 -2131
rect 129 -2199 187 -2165
rect 129 -2233 141 -2199
rect 175 -2233 187 -2199
rect 129 -2267 187 -2233
rect 129 -2301 141 -2267
rect 175 -2301 187 -2267
rect 129 -2335 187 -2301
rect 129 -2369 141 -2335
rect 175 -2369 187 -2335
rect 129 -2403 187 -2369
rect 129 -2437 141 -2403
rect 175 -2437 187 -2403
rect 129 -2471 187 -2437
rect 129 -2505 141 -2471
rect 175 -2505 187 -2471
rect 129 -2539 187 -2505
rect 129 -2573 141 -2539
rect 175 -2573 187 -2539
rect 129 -2612 187 -2573
rect 287 -1451 345 -1412
rect 287 -1485 299 -1451
rect 333 -1485 345 -1451
rect 287 -1519 345 -1485
rect 287 -1553 299 -1519
rect 333 -1553 345 -1519
rect 287 -1587 345 -1553
rect 287 -1621 299 -1587
rect 333 -1621 345 -1587
rect 287 -1655 345 -1621
rect 287 -1689 299 -1655
rect 333 -1689 345 -1655
rect 287 -1723 345 -1689
rect 287 -1757 299 -1723
rect 333 -1757 345 -1723
rect 287 -1791 345 -1757
rect 287 -1825 299 -1791
rect 333 -1825 345 -1791
rect 287 -1859 345 -1825
rect 287 -1893 299 -1859
rect 333 -1893 345 -1859
rect 287 -1927 345 -1893
rect 287 -1961 299 -1927
rect 333 -1961 345 -1927
rect 287 -1995 345 -1961
rect 287 -2029 299 -1995
rect 333 -2029 345 -1995
rect 287 -2063 345 -2029
rect 287 -2097 299 -2063
rect 333 -2097 345 -2063
rect 287 -2131 345 -2097
rect 287 -2165 299 -2131
rect 333 -2165 345 -2131
rect 287 -2199 345 -2165
rect 287 -2233 299 -2199
rect 333 -2233 345 -2199
rect 287 -2267 345 -2233
rect 287 -2301 299 -2267
rect 333 -2301 345 -2267
rect 287 -2335 345 -2301
rect 287 -2369 299 -2335
rect 333 -2369 345 -2335
rect 287 -2403 345 -2369
rect 287 -2437 299 -2403
rect 333 -2437 345 -2403
rect 287 -2471 345 -2437
rect 287 -2505 299 -2471
rect 333 -2505 345 -2471
rect 287 -2539 345 -2505
rect 287 -2573 299 -2539
rect 333 -2573 345 -2539
rect 287 -2612 345 -2573
rect 445 -1451 503 -1412
rect 445 -1485 457 -1451
rect 491 -1485 503 -1451
rect 445 -1519 503 -1485
rect 445 -1553 457 -1519
rect 491 -1553 503 -1519
rect 445 -1587 503 -1553
rect 445 -1621 457 -1587
rect 491 -1621 503 -1587
rect 445 -1655 503 -1621
rect 445 -1689 457 -1655
rect 491 -1689 503 -1655
rect 445 -1723 503 -1689
rect 445 -1757 457 -1723
rect 491 -1757 503 -1723
rect 445 -1791 503 -1757
rect 445 -1825 457 -1791
rect 491 -1825 503 -1791
rect 445 -1859 503 -1825
rect 445 -1893 457 -1859
rect 491 -1893 503 -1859
rect 445 -1927 503 -1893
rect 445 -1961 457 -1927
rect 491 -1961 503 -1927
rect 445 -1995 503 -1961
rect 445 -2029 457 -1995
rect 491 -2029 503 -1995
rect 445 -2063 503 -2029
rect 445 -2097 457 -2063
rect 491 -2097 503 -2063
rect 445 -2131 503 -2097
rect 445 -2165 457 -2131
rect 491 -2165 503 -2131
rect 445 -2199 503 -2165
rect 445 -2233 457 -2199
rect 491 -2233 503 -2199
rect 445 -2267 503 -2233
rect 445 -2301 457 -2267
rect 491 -2301 503 -2267
rect 445 -2335 503 -2301
rect 445 -2369 457 -2335
rect 491 -2369 503 -2335
rect 445 -2403 503 -2369
rect 445 -2437 457 -2403
rect 491 -2437 503 -2403
rect 445 -2471 503 -2437
rect 445 -2505 457 -2471
rect 491 -2505 503 -2471
rect 445 -2539 503 -2505
rect 445 -2573 457 -2539
rect 491 -2573 503 -2539
rect 445 -2612 503 -2573
rect 603 -1451 661 -1412
rect 603 -1485 615 -1451
rect 649 -1485 661 -1451
rect 603 -1519 661 -1485
rect 603 -1553 615 -1519
rect 649 -1553 661 -1519
rect 603 -1587 661 -1553
rect 603 -1621 615 -1587
rect 649 -1621 661 -1587
rect 603 -1655 661 -1621
rect 603 -1689 615 -1655
rect 649 -1689 661 -1655
rect 603 -1723 661 -1689
rect 603 -1757 615 -1723
rect 649 -1757 661 -1723
rect 603 -1791 661 -1757
rect 603 -1825 615 -1791
rect 649 -1825 661 -1791
rect 603 -1859 661 -1825
rect 603 -1893 615 -1859
rect 649 -1893 661 -1859
rect 603 -1927 661 -1893
rect 603 -1961 615 -1927
rect 649 -1961 661 -1927
rect 603 -1995 661 -1961
rect 603 -2029 615 -1995
rect 649 -2029 661 -1995
rect 603 -2063 661 -2029
rect 603 -2097 615 -2063
rect 649 -2097 661 -2063
rect 603 -2131 661 -2097
rect 603 -2165 615 -2131
rect 649 -2165 661 -2131
rect 603 -2199 661 -2165
rect 603 -2233 615 -2199
rect 649 -2233 661 -2199
rect 603 -2267 661 -2233
rect 603 -2301 615 -2267
rect 649 -2301 661 -2267
rect 603 -2335 661 -2301
rect 603 -2369 615 -2335
rect 649 -2369 661 -2335
rect 603 -2403 661 -2369
rect 603 -2437 615 -2403
rect 649 -2437 661 -2403
rect 603 -2471 661 -2437
rect 603 -2505 615 -2471
rect 649 -2505 661 -2471
rect 603 -2539 661 -2505
rect 603 -2573 615 -2539
rect 649 -2573 661 -2539
rect 603 -2612 661 -2573
rect 761 -1451 819 -1412
rect 761 -1485 773 -1451
rect 807 -1485 819 -1451
rect 761 -1519 819 -1485
rect 761 -1553 773 -1519
rect 807 -1553 819 -1519
rect 761 -1587 819 -1553
rect 761 -1621 773 -1587
rect 807 -1621 819 -1587
rect 761 -1655 819 -1621
rect 761 -1689 773 -1655
rect 807 -1689 819 -1655
rect 761 -1723 819 -1689
rect 761 -1757 773 -1723
rect 807 -1757 819 -1723
rect 761 -1791 819 -1757
rect 761 -1825 773 -1791
rect 807 -1825 819 -1791
rect 761 -1859 819 -1825
rect 761 -1893 773 -1859
rect 807 -1893 819 -1859
rect 761 -1927 819 -1893
rect 761 -1961 773 -1927
rect 807 -1961 819 -1927
rect 761 -1995 819 -1961
rect 761 -2029 773 -1995
rect 807 -2029 819 -1995
rect 761 -2063 819 -2029
rect 761 -2097 773 -2063
rect 807 -2097 819 -2063
rect 761 -2131 819 -2097
rect 761 -2165 773 -2131
rect 807 -2165 819 -2131
rect 761 -2199 819 -2165
rect 761 -2233 773 -2199
rect 807 -2233 819 -2199
rect 761 -2267 819 -2233
rect 761 -2301 773 -2267
rect 807 -2301 819 -2267
rect 761 -2335 819 -2301
rect 761 -2369 773 -2335
rect 807 -2369 819 -2335
rect 761 -2403 819 -2369
rect 761 -2437 773 -2403
rect 807 -2437 819 -2403
rect 761 -2471 819 -2437
rect 761 -2505 773 -2471
rect 807 -2505 819 -2471
rect 761 -2539 819 -2505
rect 761 -2573 773 -2539
rect 807 -2573 819 -2539
rect 761 -2612 819 -2573
rect 919 -1451 977 -1412
rect 919 -1485 931 -1451
rect 965 -1485 977 -1451
rect 919 -1519 977 -1485
rect 919 -1553 931 -1519
rect 965 -1553 977 -1519
rect 919 -1587 977 -1553
rect 919 -1621 931 -1587
rect 965 -1621 977 -1587
rect 919 -1655 977 -1621
rect 919 -1689 931 -1655
rect 965 -1689 977 -1655
rect 919 -1723 977 -1689
rect 919 -1757 931 -1723
rect 965 -1757 977 -1723
rect 919 -1791 977 -1757
rect 919 -1825 931 -1791
rect 965 -1825 977 -1791
rect 919 -1859 977 -1825
rect 919 -1893 931 -1859
rect 965 -1893 977 -1859
rect 919 -1927 977 -1893
rect 919 -1961 931 -1927
rect 965 -1961 977 -1927
rect 919 -1995 977 -1961
rect 919 -2029 931 -1995
rect 965 -2029 977 -1995
rect 919 -2063 977 -2029
rect 919 -2097 931 -2063
rect 965 -2097 977 -2063
rect 919 -2131 977 -2097
rect 919 -2165 931 -2131
rect 965 -2165 977 -2131
rect 919 -2199 977 -2165
rect 919 -2233 931 -2199
rect 965 -2233 977 -2199
rect 919 -2267 977 -2233
rect 919 -2301 931 -2267
rect 965 -2301 977 -2267
rect 919 -2335 977 -2301
rect 919 -2369 931 -2335
rect 965 -2369 977 -2335
rect 919 -2403 977 -2369
rect 919 -2437 931 -2403
rect 965 -2437 977 -2403
rect 919 -2471 977 -2437
rect 919 -2505 931 -2471
rect 965 -2505 977 -2471
rect 919 -2539 977 -2505
rect 919 -2573 931 -2539
rect 965 -2573 977 -2539
rect 919 -2612 977 -2573
rect 1077 -1451 1135 -1412
rect 1077 -1485 1089 -1451
rect 1123 -1485 1135 -1451
rect 1077 -1519 1135 -1485
rect 1077 -1553 1089 -1519
rect 1123 -1553 1135 -1519
rect 1077 -1587 1135 -1553
rect 1077 -1621 1089 -1587
rect 1123 -1621 1135 -1587
rect 1077 -1655 1135 -1621
rect 1077 -1689 1089 -1655
rect 1123 -1689 1135 -1655
rect 1077 -1723 1135 -1689
rect 1077 -1757 1089 -1723
rect 1123 -1757 1135 -1723
rect 1077 -1791 1135 -1757
rect 1077 -1825 1089 -1791
rect 1123 -1825 1135 -1791
rect 1077 -1859 1135 -1825
rect 1077 -1893 1089 -1859
rect 1123 -1893 1135 -1859
rect 1077 -1927 1135 -1893
rect 1077 -1961 1089 -1927
rect 1123 -1961 1135 -1927
rect 1077 -1995 1135 -1961
rect 1077 -2029 1089 -1995
rect 1123 -2029 1135 -1995
rect 1077 -2063 1135 -2029
rect 1077 -2097 1089 -2063
rect 1123 -2097 1135 -2063
rect 1077 -2131 1135 -2097
rect 1077 -2165 1089 -2131
rect 1123 -2165 1135 -2131
rect 1077 -2199 1135 -2165
rect 1077 -2233 1089 -2199
rect 1123 -2233 1135 -2199
rect 1077 -2267 1135 -2233
rect 1077 -2301 1089 -2267
rect 1123 -2301 1135 -2267
rect 1077 -2335 1135 -2301
rect 1077 -2369 1089 -2335
rect 1123 -2369 1135 -2335
rect 1077 -2403 1135 -2369
rect 1077 -2437 1089 -2403
rect 1123 -2437 1135 -2403
rect 1077 -2471 1135 -2437
rect 1077 -2505 1089 -2471
rect 1123 -2505 1135 -2471
rect 1077 -2539 1135 -2505
rect 1077 -2573 1089 -2539
rect 1123 -2573 1135 -2539
rect 1077 -2612 1135 -2573
<< pdiffc >>
rect -1123 2610 -1089 2644
rect -1123 2542 -1089 2576
rect -1123 2474 -1089 2508
rect -1123 2406 -1089 2440
rect -1123 2338 -1089 2372
rect -1123 2270 -1089 2304
rect -1123 2202 -1089 2236
rect -1123 2134 -1089 2168
rect -1123 2066 -1089 2100
rect -1123 1998 -1089 2032
rect -1123 1930 -1089 1964
rect -1123 1862 -1089 1896
rect -1123 1794 -1089 1828
rect -1123 1726 -1089 1760
rect -1123 1658 -1089 1692
rect -1123 1590 -1089 1624
rect -1123 1522 -1089 1556
rect -965 2610 -931 2644
rect -965 2542 -931 2576
rect -965 2474 -931 2508
rect -965 2406 -931 2440
rect -965 2338 -931 2372
rect -965 2270 -931 2304
rect -965 2202 -931 2236
rect -965 2134 -931 2168
rect -965 2066 -931 2100
rect -965 1998 -931 2032
rect -965 1930 -931 1964
rect -965 1862 -931 1896
rect -965 1794 -931 1828
rect -965 1726 -931 1760
rect -965 1658 -931 1692
rect -965 1590 -931 1624
rect -965 1522 -931 1556
rect -807 2610 -773 2644
rect -807 2542 -773 2576
rect -807 2474 -773 2508
rect -807 2406 -773 2440
rect -807 2338 -773 2372
rect -807 2270 -773 2304
rect -807 2202 -773 2236
rect -807 2134 -773 2168
rect -807 2066 -773 2100
rect -807 1998 -773 2032
rect -807 1930 -773 1964
rect -807 1862 -773 1896
rect -807 1794 -773 1828
rect -807 1726 -773 1760
rect -807 1658 -773 1692
rect -807 1590 -773 1624
rect -807 1522 -773 1556
rect -649 2610 -615 2644
rect -649 2542 -615 2576
rect -649 2474 -615 2508
rect -649 2406 -615 2440
rect -649 2338 -615 2372
rect -649 2270 -615 2304
rect -649 2202 -615 2236
rect -649 2134 -615 2168
rect -649 2066 -615 2100
rect -649 1998 -615 2032
rect -649 1930 -615 1964
rect -649 1862 -615 1896
rect -649 1794 -615 1828
rect -649 1726 -615 1760
rect -649 1658 -615 1692
rect -649 1590 -615 1624
rect -649 1522 -615 1556
rect -491 2610 -457 2644
rect -491 2542 -457 2576
rect -491 2474 -457 2508
rect -491 2406 -457 2440
rect -491 2338 -457 2372
rect -491 2270 -457 2304
rect -491 2202 -457 2236
rect -491 2134 -457 2168
rect -491 2066 -457 2100
rect -491 1998 -457 2032
rect -491 1930 -457 1964
rect -491 1862 -457 1896
rect -491 1794 -457 1828
rect -491 1726 -457 1760
rect -491 1658 -457 1692
rect -491 1590 -457 1624
rect -491 1522 -457 1556
rect -333 2610 -299 2644
rect -333 2542 -299 2576
rect -333 2474 -299 2508
rect -333 2406 -299 2440
rect -333 2338 -299 2372
rect -333 2270 -299 2304
rect -333 2202 -299 2236
rect -333 2134 -299 2168
rect -333 2066 -299 2100
rect -333 1998 -299 2032
rect -333 1930 -299 1964
rect -333 1862 -299 1896
rect -333 1794 -299 1828
rect -333 1726 -299 1760
rect -333 1658 -299 1692
rect -333 1590 -299 1624
rect -333 1522 -299 1556
rect -175 2610 -141 2644
rect -175 2542 -141 2576
rect -175 2474 -141 2508
rect -175 2406 -141 2440
rect -175 2338 -141 2372
rect -175 2270 -141 2304
rect -175 2202 -141 2236
rect -175 2134 -141 2168
rect -175 2066 -141 2100
rect -175 1998 -141 2032
rect -175 1930 -141 1964
rect -175 1862 -141 1896
rect -175 1794 -141 1828
rect -175 1726 -141 1760
rect -175 1658 -141 1692
rect -175 1590 -141 1624
rect -175 1522 -141 1556
rect -17 2610 17 2644
rect -17 2542 17 2576
rect -17 2474 17 2508
rect -17 2406 17 2440
rect -17 2338 17 2372
rect -17 2270 17 2304
rect -17 2202 17 2236
rect -17 2134 17 2168
rect -17 2066 17 2100
rect -17 1998 17 2032
rect -17 1930 17 1964
rect -17 1862 17 1896
rect -17 1794 17 1828
rect -17 1726 17 1760
rect -17 1658 17 1692
rect -17 1590 17 1624
rect -17 1522 17 1556
rect 141 2610 175 2644
rect 141 2542 175 2576
rect 141 2474 175 2508
rect 141 2406 175 2440
rect 141 2338 175 2372
rect 141 2270 175 2304
rect 141 2202 175 2236
rect 141 2134 175 2168
rect 141 2066 175 2100
rect 141 1998 175 2032
rect 141 1930 175 1964
rect 141 1862 175 1896
rect 141 1794 175 1828
rect 141 1726 175 1760
rect 141 1658 175 1692
rect 141 1590 175 1624
rect 141 1522 175 1556
rect 299 2610 333 2644
rect 299 2542 333 2576
rect 299 2474 333 2508
rect 299 2406 333 2440
rect 299 2338 333 2372
rect 299 2270 333 2304
rect 299 2202 333 2236
rect 299 2134 333 2168
rect 299 2066 333 2100
rect 299 1998 333 2032
rect 299 1930 333 1964
rect 299 1862 333 1896
rect 299 1794 333 1828
rect 299 1726 333 1760
rect 299 1658 333 1692
rect 299 1590 333 1624
rect 299 1522 333 1556
rect 457 2610 491 2644
rect 457 2542 491 2576
rect 457 2474 491 2508
rect 457 2406 491 2440
rect 457 2338 491 2372
rect 457 2270 491 2304
rect 457 2202 491 2236
rect 457 2134 491 2168
rect 457 2066 491 2100
rect 457 1998 491 2032
rect 457 1930 491 1964
rect 457 1862 491 1896
rect 457 1794 491 1828
rect 457 1726 491 1760
rect 457 1658 491 1692
rect 457 1590 491 1624
rect 457 1522 491 1556
rect 615 2610 649 2644
rect 615 2542 649 2576
rect 615 2474 649 2508
rect 615 2406 649 2440
rect 615 2338 649 2372
rect 615 2270 649 2304
rect 615 2202 649 2236
rect 615 2134 649 2168
rect 615 2066 649 2100
rect 615 1998 649 2032
rect 615 1930 649 1964
rect 615 1862 649 1896
rect 615 1794 649 1828
rect 615 1726 649 1760
rect 615 1658 649 1692
rect 615 1590 649 1624
rect 615 1522 649 1556
rect 773 2610 807 2644
rect 773 2542 807 2576
rect 773 2474 807 2508
rect 773 2406 807 2440
rect 773 2338 807 2372
rect 773 2270 807 2304
rect 773 2202 807 2236
rect 773 2134 807 2168
rect 773 2066 807 2100
rect 773 1998 807 2032
rect 773 1930 807 1964
rect 773 1862 807 1896
rect 773 1794 807 1828
rect 773 1726 807 1760
rect 773 1658 807 1692
rect 773 1590 807 1624
rect 773 1522 807 1556
rect 931 2610 965 2644
rect 931 2542 965 2576
rect 931 2474 965 2508
rect 931 2406 965 2440
rect 931 2338 965 2372
rect 931 2270 965 2304
rect 931 2202 965 2236
rect 931 2134 965 2168
rect 931 2066 965 2100
rect 931 1998 965 2032
rect 931 1930 965 1964
rect 931 1862 965 1896
rect 931 1794 965 1828
rect 931 1726 965 1760
rect 931 1658 965 1692
rect 931 1590 965 1624
rect 931 1522 965 1556
rect 1089 2610 1123 2644
rect 1089 2542 1123 2576
rect 1089 2474 1123 2508
rect 1089 2406 1123 2440
rect 1089 2338 1123 2372
rect 1089 2270 1123 2304
rect 1089 2202 1123 2236
rect 1089 2134 1123 2168
rect 1089 2066 1123 2100
rect 1089 1998 1123 2032
rect 1089 1930 1123 1964
rect 1089 1862 1123 1896
rect 1089 1794 1123 1828
rect 1089 1726 1123 1760
rect 1089 1658 1123 1692
rect 1089 1590 1123 1624
rect 1089 1522 1123 1556
rect -1123 1245 -1089 1279
rect -1123 1177 -1089 1211
rect -1123 1109 -1089 1143
rect -1123 1041 -1089 1075
rect -1123 973 -1089 1007
rect -1123 905 -1089 939
rect -1123 837 -1089 871
rect -1123 769 -1089 803
rect -1123 701 -1089 735
rect -1123 633 -1089 667
rect -1123 565 -1089 599
rect -1123 497 -1089 531
rect -1123 429 -1089 463
rect -1123 361 -1089 395
rect -1123 293 -1089 327
rect -1123 225 -1089 259
rect -1123 157 -1089 191
rect -965 1245 -931 1279
rect -965 1177 -931 1211
rect -965 1109 -931 1143
rect -965 1041 -931 1075
rect -965 973 -931 1007
rect -965 905 -931 939
rect -965 837 -931 871
rect -965 769 -931 803
rect -965 701 -931 735
rect -965 633 -931 667
rect -965 565 -931 599
rect -965 497 -931 531
rect -965 429 -931 463
rect -965 361 -931 395
rect -965 293 -931 327
rect -965 225 -931 259
rect -965 157 -931 191
rect -807 1245 -773 1279
rect -807 1177 -773 1211
rect -807 1109 -773 1143
rect -807 1041 -773 1075
rect -807 973 -773 1007
rect -807 905 -773 939
rect -807 837 -773 871
rect -807 769 -773 803
rect -807 701 -773 735
rect -807 633 -773 667
rect -807 565 -773 599
rect -807 497 -773 531
rect -807 429 -773 463
rect -807 361 -773 395
rect -807 293 -773 327
rect -807 225 -773 259
rect -807 157 -773 191
rect -649 1245 -615 1279
rect -649 1177 -615 1211
rect -649 1109 -615 1143
rect -649 1041 -615 1075
rect -649 973 -615 1007
rect -649 905 -615 939
rect -649 837 -615 871
rect -649 769 -615 803
rect -649 701 -615 735
rect -649 633 -615 667
rect -649 565 -615 599
rect -649 497 -615 531
rect -649 429 -615 463
rect -649 361 -615 395
rect -649 293 -615 327
rect -649 225 -615 259
rect -649 157 -615 191
rect -491 1245 -457 1279
rect -491 1177 -457 1211
rect -491 1109 -457 1143
rect -491 1041 -457 1075
rect -491 973 -457 1007
rect -491 905 -457 939
rect -491 837 -457 871
rect -491 769 -457 803
rect -491 701 -457 735
rect -491 633 -457 667
rect -491 565 -457 599
rect -491 497 -457 531
rect -491 429 -457 463
rect -491 361 -457 395
rect -491 293 -457 327
rect -491 225 -457 259
rect -491 157 -457 191
rect -333 1245 -299 1279
rect -333 1177 -299 1211
rect -333 1109 -299 1143
rect -333 1041 -299 1075
rect -333 973 -299 1007
rect -333 905 -299 939
rect -333 837 -299 871
rect -333 769 -299 803
rect -333 701 -299 735
rect -333 633 -299 667
rect -333 565 -299 599
rect -333 497 -299 531
rect -333 429 -299 463
rect -333 361 -299 395
rect -333 293 -299 327
rect -333 225 -299 259
rect -333 157 -299 191
rect -175 1245 -141 1279
rect -175 1177 -141 1211
rect -175 1109 -141 1143
rect -175 1041 -141 1075
rect -175 973 -141 1007
rect -175 905 -141 939
rect -175 837 -141 871
rect -175 769 -141 803
rect -175 701 -141 735
rect -175 633 -141 667
rect -175 565 -141 599
rect -175 497 -141 531
rect -175 429 -141 463
rect -175 361 -141 395
rect -175 293 -141 327
rect -175 225 -141 259
rect -175 157 -141 191
rect -17 1245 17 1279
rect -17 1177 17 1211
rect -17 1109 17 1143
rect -17 1041 17 1075
rect -17 973 17 1007
rect -17 905 17 939
rect -17 837 17 871
rect -17 769 17 803
rect -17 701 17 735
rect -17 633 17 667
rect -17 565 17 599
rect -17 497 17 531
rect -17 429 17 463
rect -17 361 17 395
rect -17 293 17 327
rect -17 225 17 259
rect -17 157 17 191
rect 141 1245 175 1279
rect 141 1177 175 1211
rect 141 1109 175 1143
rect 141 1041 175 1075
rect 141 973 175 1007
rect 141 905 175 939
rect 141 837 175 871
rect 141 769 175 803
rect 141 701 175 735
rect 141 633 175 667
rect 141 565 175 599
rect 141 497 175 531
rect 141 429 175 463
rect 141 361 175 395
rect 141 293 175 327
rect 141 225 175 259
rect 141 157 175 191
rect 299 1245 333 1279
rect 299 1177 333 1211
rect 299 1109 333 1143
rect 299 1041 333 1075
rect 299 973 333 1007
rect 299 905 333 939
rect 299 837 333 871
rect 299 769 333 803
rect 299 701 333 735
rect 299 633 333 667
rect 299 565 333 599
rect 299 497 333 531
rect 299 429 333 463
rect 299 361 333 395
rect 299 293 333 327
rect 299 225 333 259
rect 299 157 333 191
rect 457 1245 491 1279
rect 457 1177 491 1211
rect 457 1109 491 1143
rect 457 1041 491 1075
rect 457 973 491 1007
rect 457 905 491 939
rect 457 837 491 871
rect 457 769 491 803
rect 457 701 491 735
rect 457 633 491 667
rect 457 565 491 599
rect 457 497 491 531
rect 457 429 491 463
rect 457 361 491 395
rect 457 293 491 327
rect 457 225 491 259
rect 457 157 491 191
rect 615 1245 649 1279
rect 615 1177 649 1211
rect 615 1109 649 1143
rect 615 1041 649 1075
rect 615 973 649 1007
rect 615 905 649 939
rect 615 837 649 871
rect 615 769 649 803
rect 615 701 649 735
rect 615 633 649 667
rect 615 565 649 599
rect 615 497 649 531
rect 615 429 649 463
rect 615 361 649 395
rect 615 293 649 327
rect 615 225 649 259
rect 615 157 649 191
rect 773 1245 807 1279
rect 773 1177 807 1211
rect 773 1109 807 1143
rect 773 1041 807 1075
rect 773 973 807 1007
rect 773 905 807 939
rect 773 837 807 871
rect 773 769 807 803
rect 773 701 807 735
rect 773 633 807 667
rect 773 565 807 599
rect 773 497 807 531
rect 773 429 807 463
rect 773 361 807 395
rect 773 293 807 327
rect 773 225 807 259
rect 773 157 807 191
rect 931 1245 965 1279
rect 931 1177 965 1211
rect 931 1109 965 1143
rect 931 1041 965 1075
rect 931 973 965 1007
rect 931 905 965 939
rect 931 837 965 871
rect 931 769 965 803
rect 931 701 965 735
rect 931 633 965 667
rect 931 565 965 599
rect 931 497 965 531
rect 931 429 965 463
rect 931 361 965 395
rect 931 293 965 327
rect 931 225 965 259
rect 931 157 965 191
rect 1089 1245 1123 1279
rect 1089 1177 1123 1211
rect 1089 1109 1123 1143
rect 1089 1041 1123 1075
rect 1089 973 1123 1007
rect 1089 905 1123 939
rect 1089 837 1123 871
rect 1089 769 1123 803
rect 1089 701 1123 735
rect 1089 633 1123 667
rect 1089 565 1123 599
rect 1089 497 1123 531
rect 1089 429 1123 463
rect 1089 361 1123 395
rect 1089 293 1123 327
rect 1089 225 1123 259
rect 1089 157 1123 191
rect -1123 -120 -1089 -86
rect -1123 -188 -1089 -154
rect -1123 -256 -1089 -222
rect -1123 -324 -1089 -290
rect -1123 -392 -1089 -358
rect -1123 -460 -1089 -426
rect -1123 -528 -1089 -494
rect -1123 -596 -1089 -562
rect -1123 -664 -1089 -630
rect -1123 -732 -1089 -698
rect -1123 -800 -1089 -766
rect -1123 -868 -1089 -834
rect -1123 -936 -1089 -902
rect -1123 -1004 -1089 -970
rect -1123 -1072 -1089 -1038
rect -1123 -1140 -1089 -1106
rect -1123 -1208 -1089 -1174
rect -965 -120 -931 -86
rect -965 -188 -931 -154
rect -965 -256 -931 -222
rect -965 -324 -931 -290
rect -965 -392 -931 -358
rect -965 -460 -931 -426
rect -965 -528 -931 -494
rect -965 -596 -931 -562
rect -965 -664 -931 -630
rect -965 -732 -931 -698
rect -965 -800 -931 -766
rect -965 -868 -931 -834
rect -965 -936 -931 -902
rect -965 -1004 -931 -970
rect -965 -1072 -931 -1038
rect -965 -1140 -931 -1106
rect -965 -1208 -931 -1174
rect -807 -120 -773 -86
rect -807 -188 -773 -154
rect -807 -256 -773 -222
rect -807 -324 -773 -290
rect -807 -392 -773 -358
rect -807 -460 -773 -426
rect -807 -528 -773 -494
rect -807 -596 -773 -562
rect -807 -664 -773 -630
rect -807 -732 -773 -698
rect -807 -800 -773 -766
rect -807 -868 -773 -834
rect -807 -936 -773 -902
rect -807 -1004 -773 -970
rect -807 -1072 -773 -1038
rect -807 -1140 -773 -1106
rect -807 -1208 -773 -1174
rect -649 -120 -615 -86
rect -649 -188 -615 -154
rect -649 -256 -615 -222
rect -649 -324 -615 -290
rect -649 -392 -615 -358
rect -649 -460 -615 -426
rect -649 -528 -615 -494
rect -649 -596 -615 -562
rect -649 -664 -615 -630
rect -649 -732 -615 -698
rect -649 -800 -615 -766
rect -649 -868 -615 -834
rect -649 -936 -615 -902
rect -649 -1004 -615 -970
rect -649 -1072 -615 -1038
rect -649 -1140 -615 -1106
rect -649 -1208 -615 -1174
rect -491 -120 -457 -86
rect -491 -188 -457 -154
rect -491 -256 -457 -222
rect -491 -324 -457 -290
rect -491 -392 -457 -358
rect -491 -460 -457 -426
rect -491 -528 -457 -494
rect -491 -596 -457 -562
rect -491 -664 -457 -630
rect -491 -732 -457 -698
rect -491 -800 -457 -766
rect -491 -868 -457 -834
rect -491 -936 -457 -902
rect -491 -1004 -457 -970
rect -491 -1072 -457 -1038
rect -491 -1140 -457 -1106
rect -491 -1208 -457 -1174
rect -333 -120 -299 -86
rect -333 -188 -299 -154
rect -333 -256 -299 -222
rect -333 -324 -299 -290
rect -333 -392 -299 -358
rect -333 -460 -299 -426
rect -333 -528 -299 -494
rect -333 -596 -299 -562
rect -333 -664 -299 -630
rect -333 -732 -299 -698
rect -333 -800 -299 -766
rect -333 -868 -299 -834
rect -333 -936 -299 -902
rect -333 -1004 -299 -970
rect -333 -1072 -299 -1038
rect -333 -1140 -299 -1106
rect -333 -1208 -299 -1174
rect -175 -120 -141 -86
rect -175 -188 -141 -154
rect -175 -256 -141 -222
rect -175 -324 -141 -290
rect -175 -392 -141 -358
rect -175 -460 -141 -426
rect -175 -528 -141 -494
rect -175 -596 -141 -562
rect -175 -664 -141 -630
rect -175 -732 -141 -698
rect -175 -800 -141 -766
rect -175 -868 -141 -834
rect -175 -936 -141 -902
rect -175 -1004 -141 -970
rect -175 -1072 -141 -1038
rect -175 -1140 -141 -1106
rect -175 -1208 -141 -1174
rect -17 -120 17 -86
rect -17 -188 17 -154
rect -17 -256 17 -222
rect -17 -324 17 -290
rect -17 -392 17 -358
rect -17 -460 17 -426
rect -17 -528 17 -494
rect -17 -596 17 -562
rect -17 -664 17 -630
rect -17 -732 17 -698
rect -17 -800 17 -766
rect -17 -868 17 -834
rect -17 -936 17 -902
rect -17 -1004 17 -970
rect -17 -1072 17 -1038
rect -17 -1140 17 -1106
rect -17 -1208 17 -1174
rect 141 -120 175 -86
rect 141 -188 175 -154
rect 141 -256 175 -222
rect 141 -324 175 -290
rect 141 -392 175 -358
rect 141 -460 175 -426
rect 141 -528 175 -494
rect 141 -596 175 -562
rect 141 -664 175 -630
rect 141 -732 175 -698
rect 141 -800 175 -766
rect 141 -868 175 -834
rect 141 -936 175 -902
rect 141 -1004 175 -970
rect 141 -1072 175 -1038
rect 141 -1140 175 -1106
rect 141 -1208 175 -1174
rect 299 -120 333 -86
rect 299 -188 333 -154
rect 299 -256 333 -222
rect 299 -324 333 -290
rect 299 -392 333 -358
rect 299 -460 333 -426
rect 299 -528 333 -494
rect 299 -596 333 -562
rect 299 -664 333 -630
rect 299 -732 333 -698
rect 299 -800 333 -766
rect 299 -868 333 -834
rect 299 -936 333 -902
rect 299 -1004 333 -970
rect 299 -1072 333 -1038
rect 299 -1140 333 -1106
rect 299 -1208 333 -1174
rect 457 -120 491 -86
rect 457 -188 491 -154
rect 457 -256 491 -222
rect 457 -324 491 -290
rect 457 -392 491 -358
rect 457 -460 491 -426
rect 457 -528 491 -494
rect 457 -596 491 -562
rect 457 -664 491 -630
rect 457 -732 491 -698
rect 457 -800 491 -766
rect 457 -868 491 -834
rect 457 -936 491 -902
rect 457 -1004 491 -970
rect 457 -1072 491 -1038
rect 457 -1140 491 -1106
rect 457 -1208 491 -1174
rect 615 -120 649 -86
rect 615 -188 649 -154
rect 615 -256 649 -222
rect 615 -324 649 -290
rect 615 -392 649 -358
rect 615 -460 649 -426
rect 615 -528 649 -494
rect 615 -596 649 -562
rect 615 -664 649 -630
rect 615 -732 649 -698
rect 615 -800 649 -766
rect 615 -868 649 -834
rect 615 -936 649 -902
rect 615 -1004 649 -970
rect 615 -1072 649 -1038
rect 615 -1140 649 -1106
rect 615 -1208 649 -1174
rect 773 -120 807 -86
rect 773 -188 807 -154
rect 773 -256 807 -222
rect 773 -324 807 -290
rect 773 -392 807 -358
rect 773 -460 807 -426
rect 773 -528 807 -494
rect 773 -596 807 -562
rect 773 -664 807 -630
rect 773 -732 807 -698
rect 773 -800 807 -766
rect 773 -868 807 -834
rect 773 -936 807 -902
rect 773 -1004 807 -970
rect 773 -1072 807 -1038
rect 773 -1140 807 -1106
rect 773 -1208 807 -1174
rect 931 -120 965 -86
rect 931 -188 965 -154
rect 931 -256 965 -222
rect 931 -324 965 -290
rect 931 -392 965 -358
rect 931 -460 965 -426
rect 931 -528 965 -494
rect 931 -596 965 -562
rect 931 -664 965 -630
rect 931 -732 965 -698
rect 931 -800 965 -766
rect 931 -868 965 -834
rect 931 -936 965 -902
rect 931 -1004 965 -970
rect 931 -1072 965 -1038
rect 931 -1140 965 -1106
rect 931 -1208 965 -1174
rect 1089 -120 1123 -86
rect 1089 -188 1123 -154
rect 1089 -256 1123 -222
rect 1089 -324 1123 -290
rect 1089 -392 1123 -358
rect 1089 -460 1123 -426
rect 1089 -528 1123 -494
rect 1089 -596 1123 -562
rect 1089 -664 1123 -630
rect 1089 -732 1123 -698
rect 1089 -800 1123 -766
rect 1089 -868 1123 -834
rect 1089 -936 1123 -902
rect 1089 -1004 1123 -970
rect 1089 -1072 1123 -1038
rect 1089 -1140 1123 -1106
rect 1089 -1208 1123 -1174
rect -1123 -1485 -1089 -1451
rect -1123 -1553 -1089 -1519
rect -1123 -1621 -1089 -1587
rect -1123 -1689 -1089 -1655
rect -1123 -1757 -1089 -1723
rect -1123 -1825 -1089 -1791
rect -1123 -1893 -1089 -1859
rect -1123 -1961 -1089 -1927
rect -1123 -2029 -1089 -1995
rect -1123 -2097 -1089 -2063
rect -1123 -2165 -1089 -2131
rect -1123 -2233 -1089 -2199
rect -1123 -2301 -1089 -2267
rect -1123 -2369 -1089 -2335
rect -1123 -2437 -1089 -2403
rect -1123 -2505 -1089 -2471
rect -1123 -2573 -1089 -2539
rect -965 -1485 -931 -1451
rect -965 -1553 -931 -1519
rect -965 -1621 -931 -1587
rect -965 -1689 -931 -1655
rect -965 -1757 -931 -1723
rect -965 -1825 -931 -1791
rect -965 -1893 -931 -1859
rect -965 -1961 -931 -1927
rect -965 -2029 -931 -1995
rect -965 -2097 -931 -2063
rect -965 -2165 -931 -2131
rect -965 -2233 -931 -2199
rect -965 -2301 -931 -2267
rect -965 -2369 -931 -2335
rect -965 -2437 -931 -2403
rect -965 -2505 -931 -2471
rect -965 -2573 -931 -2539
rect -807 -1485 -773 -1451
rect -807 -1553 -773 -1519
rect -807 -1621 -773 -1587
rect -807 -1689 -773 -1655
rect -807 -1757 -773 -1723
rect -807 -1825 -773 -1791
rect -807 -1893 -773 -1859
rect -807 -1961 -773 -1927
rect -807 -2029 -773 -1995
rect -807 -2097 -773 -2063
rect -807 -2165 -773 -2131
rect -807 -2233 -773 -2199
rect -807 -2301 -773 -2267
rect -807 -2369 -773 -2335
rect -807 -2437 -773 -2403
rect -807 -2505 -773 -2471
rect -807 -2573 -773 -2539
rect -649 -1485 -615 -1451
rect -649 -1553 -615 -1519
rect -649 -1621 -615 -1587
rect -649 -1689 -615 -1655
rect -649 -1757 -615 -1723
rect -649 -1825 -615 -1791
rect -649 -1893 -615 -1859
rect -649 -1961 -615 -1927
rect -649 -2029 -615 -1995
rect -649 -2097 -615 -2063
rect -649 -2165 -615 -2131
rect -649 -2233 -615 -2199
rect -649 -2301 -615 -2267
rect -649 -2369 -615 -2335
rect -649 -2437 -615 -2403
rect -649 -2505 -615 -2471
rect -649 -2573 -615 -2539
rect -491 -1485 -457 -1451
rect -491 -1553 -457 -1519
rect -491 -1621 -457 -1587
rect -491 -1689 -457 -1655
rect -491 -1757 -457 -1723
rect -491 -1825 -457 -1791
rect -491 -1893 -457 -1859
rect -491 -1961 -457 -1927
rect -491 -2029 -457 -1995
rect -491 -2097 -457 -2063
rect -491 -2165 -457 -2131
rect -491 -2233 -457 -2199
rect -491 -2301 -457 -2267
rect -491 -2369 -457 -2335
rect -491 -2437 -457 -2403
rect -491 -2505 -457 -2471
rect -491 -2573 -457 -2539
rect -333 -1485 -299 -1451
rect -333 -1553 -299 -1519
rect -333 -1621 -299 -1587
rect -333 -1689 -299 -1655
rect -333 -1757 -299 -1723
rect -333 -1825 -299 -1791
rect -333 -1893 -299 -1859
rect -333 -1961 -299 -1927
rect -333 -2029 -299 -1995
rect -333 -2097 -299 -2063
rect -333 -2165 -299 -2131
rect -333 -2233 -299 -2199
rect -333 -2301 -299 -2267
rect -333 -2369 -299 -2335
rect -333 -2437 -299 -2403
rect -333 -2505 -299 -2471
rect -333 -2573 -299 -2539
rect -175 -1485 -141 -1451
rect -175 -1553 -141 -1519
rect -175 -1621 -141 -1587
rect -175 -1689 -141 -1655
rect -175 -1757 -141 -1723
rect -175 -1825 -141 -1791
rect -175 -1893 -141 -1859
rect -175 -1961 -141 -1927
rect -175 -2029 -141 -1995
rect -175 -2097 -141 -2063
rect -175 -2165 -141 -2131
rect -175 -2233 -141 -2199
rect -175 -2301 -141 -2267
rect -175 -2369 -141 -2335
rect -175 -2437 -141 -2403
rect -175 -2505 -141 -2471
rect -175 -2573 -141 -2539
rect -17 -1485 17 -1451
rect -17 -1553 17 -1519
rect -17 -1621 17 -1587
rect -17 -1689 17 -1655
rect -17 -1757 17 -1723
rect -17 -1825 17 -1791
rect -17 -1893 17 -1859
rect -17 -1961 17 -1927
rect -17 -2029 17 -1995
rect -17 -2097 17 -2063
rect -17 -2165 17 -2131
rect -17 -2233 17 -2199
rect -17 -2301 17 -2267
rect -17 -2369 17 -2335
rect -17 -2437 17 -2403
rect -17 -2505 17 -2471
rect -17 -2573 17 -2539
rect 141 -1485 175 -1451
rect 141 -1553 175 -1519
rect 141 -1621 175 -1587
rect 141 -1689 175 -1655
rect 141 -1757 175 -1723
rect 141 -1825 175 -1791
rect 141 -1893 175 -1859
rect 141 -1961 175 -1927
rect 141 -2029 175 -1995
rect 141 -2097 175 -2063
rect 141 -2165 175 -2131
rect 141 -2233 175 -2199
rect 141 -2301 175 -2267
rect 141 -2369 175 -2335
rect 141 -2437 175 -2403
rect 141 -2505 175 -2471
rect 141 -2573 175 -2539
rect 299 -1485 333 -1451
rect 299 -1553 333 -1519
rect 299 -1621 333 -1587
rect 299 -1689 333 -1655
rect 299 -1757 333 -1723
rect 299 -1825 333 -1791
rect 299 -1893 333 -1859
rect 299 -1961 333 -1927
rect 299 -2029 333 -1995
rect 299 -2097 333 -2063
rect 299 -2165 333 -2131
rect 299 -2233 333 -2199
rect 299 -2301 333 -2267
rect 299 -2369 333 -2335
rect 299 -2437 333 -2403
rect 299 -2505 333 -2471
rect 299 -2573 333 -2539
rect 457 -1485 491 -1451
rect 457 -1553 491 -1519
rect 457 -1621 491 -1587
rect 457 -1689 491 -1655
rect 457 -1757 491 -1723
rect 457 -1825 491 -1791
rect 457 -1893 491 -1859
rect 457 -1961 491 -1927
rect 457 -2029 491 -1995
rect 457 -2097 491 -2063
rect 457 -2165 491 -2131
rect 457 -2233 491 -2199
rect 457 -2301 491 -2267
rect 457 -2369 491 -2335
rect 457 -2437 491 -2403
rect 457 -2505 491 -2471
rect 457 -2573 491 -2539
rect 615 -1485 649 -1451
rect 615 -1553 649 -1519
rect 615 -1621 649 -1587
rect 615 -1689 649 -1655
rect 615 -1757 649 -1723
rect 615 -1825 649 -1791
rect 615 -1893 649 -1859
rect 615 -1961 649 -1927
rect 615 -2029 649 -1995
rect 615 -2097 649 -2063
rect 615 -2165 649 -2131
rect 615 -2233 649 -2199
rect 615 -2301 649 -2267
rect 615 -2369 649 -2335
rect 615 -2437 649 -2403
rect 615 -2505 649 -2471
rect 615 -2573 649 -2539
rect 773 -1485 807 -1451
rect 773 -1553 807 -1519
rect 773 -1621 807 -1587
rect 773 -1689 807 -1655
rect 773 -1757 807 -1723
rect 773 -1825 807 -1791
rect 773 -1893 807 -1859
rect 773 -1961 807 -1927
rect 773 -2029 807 -1995
rect 773 -2097 807 -2063
rect 773 -2165 807 -2131
rect 773 -2233 807 -2199
rect 773 -2301 807 -2267
rect 773 -2369 807 -2335
rect 773 -2437 807 -2403
rect 773 -2505 807 -2471
rect 773 -2573 807 -2539
rect 931 -1485 965 -1451
rect 931 -1553 965 -1519
rect 931 -1621 965 -1587
rect 931 -1689 965 -1655
rect 931 -1757 965 -1723
rect 931 -1825 965 -1791
rect 931 -1893 965 -1859
rect 931 -1961 965 -1927
rect 931 -2029 965 -1995
rect 931 -2097 965 -2063
rect 931 -2165 965 -2131
rect 931 -2233 965 -2199
rect 931 -2301 965 -2267
rect 931 -2369 965 -2335
rect 931 -2437 965 -2403
rect 931 -2505 965 -2471
rect 931 -2573 965 -2539
rect 1089 -1485 1123 -1451
rect 1089 -1553 1123 -1519
rect 1089 -1621 1123 -1587
rect 1089 -1689 1123 -1655
rect 1089 -1757 1123 -1723
rect 1089 -1825 1123 -1791
rect 1089 -1893 1123 -1859
rect 1089 -1961 1123 -1927
rect 1089 -2029 1123 -1995
rect 1089 -2097 1123 -2063
rect 1089 -2165 1123 -2131
rect 1089 -2233 1123 -2199
rect 1089 -2301 1123 -2267
rect 1089 -2369 1123 -2335
rect 1089 -2437 1123 -2403
rect 1089 -2505 1123 -2471
rect 1089 -2573 1123 -2539
<< nsubdiff >>
rect -1237 2761 -1139 2795
rect -1105 2761 -1071 2795
rect -1037 2761 -1003 2795
rect -969 2761 -935 2795
rect -901 2761 -867 2795
rect -833 2761 -799 2795
rect -765 2761 -731 2795
rect -697 2761 -663 2795
rect -629 2761 -595 2795
rect -561 2761 -527 2795
rect -493 2761 -459 2795
rect -425 2761 -391 2795
rect -357 2761 -323 2795
rect -289 2761 -255 2795
rect -221 2761 -187 2795
rect -153 2761 -119 2795
rect -85 2761 -51 2795
rect -17 2761 17 2795
rect 51 2761 85 2795
rect 119 2761 153 2795
rect 187 2761 221 2795
rect 255 2761 289 2795
rect 323 2761 357 2795
rect 391 2761 425 2795
rect 459 2761 493 2795
rect 527 2761 561 2795
rect 595 2761 629 2795
rect 663 2761 697 2795
rect 731 2761 765 2795
rect 799 2761 833 2795
rect 867 2761 901 2795
rect 935 2761 969 2795
rect 1003 2761 1037 2795
rect 1071 2761 1105 2795
rect 1139 2761 1237 2795
rect -1237 2669 -1203 2761
rect -1237 2601 -1203 2635
rect -1237 2533 -1203 2567
rect -1237 2465 -1203 2499
rect -1237 2397 -1203 2431
rect -1237 2329 -1203 2363
rect -1237 2261 -1203 2295
rect -1237 2193 -1203 2227
rect -1237 2125 -1203 2159
rect -1237 2057 -1203 2091
rect -1237 1989 -1203 2023
rect -1237 1921 -1203 1955
rect -1237 1853 -1203 1887
rect -1237 1785 -1203 1819
rect -1237 1717 -1203 1751
rect -1237 1649 -1203 1683
rect -1237 1581 -1203 1615
rect -1237 1513 -1203 1547
rect 1203 2669 1237 2761
rect 1203 2601 1237 2635
rect 1203 2533 1237 2567
rect 1203 2465 1237 2499
rect 1203 2397 1237 2431
rect 1203 2329 1237 2363
rect 1203 2261 1237 2295
rect 1203 2193 1237 2227
rect 1203 2125 1237 2159
rect 1203 2057 1237 2091
rect 1203 1989 1237 2023
rect 1203 1921 1237 1955
rect 1203 1853 1237 1887
rect 1203 1785 1237 1819
rect 1203 1717 1237 1751
rect 1203 1649 1237 1683
rect 1203 1581 1237 1615
rect 1203 1513 1237 1547
rect -1237 1445 -1203 1479
rect -1237 1377 -1203 1411
rect 1203 1445 1237 1479
rect 1203 1377 1237 1411
rect -1237 1309 -1203 1343
rect -1237 1241 -1203 1275
rect -1237 1173 -1203 1207
rect -1237 1105 -1203 1139
rect -1237 1037 -1203 1071
rect -1237 969 -1203 1003
rect -1237 901 -1203 935
rect -1237 833 -1203 867
rect -1237 765 -1203 799
rect -1237 697 -1203 731
rect -1237 629 -1203 663
rect -1237 561 -1203 595
rect -1237 493 -1203 527
rect -1237 425 -1203 459
rect -1237 357 -1203 391
rect -1237 289 -1203 323
rect -1237 221 -1203 255
rect -1237 153 -1203 187
rect -1237 85 -1203 119
rect 1203 1309 1237 1343
rect 1203 1241 1237 1275
rect 1203 1173 1237 1207
rect 1203 1105 1237 1139
rect 1203 1037 1237 1071
rect 1203 969 1237 1003
rect 1203 901 1237 935
rect 1203 833 1237 867
rect 1203 765 1237 799
rect 1203 697 1237 731
rect 1203 629 1237 663
rect 1203 561 1237 595
rect 1203 493 1237 527
rect 1203 425 1237 459
rect 1203 357 1237 391
rect 1203 289 1237 323
rect 1203 221 1237 255
rect 1203 153 1237 187
rect -1237 17 -1203 51
rect 1203 85 1237 119
rect -1237 -51 -1203 -17
rect 1203 17 1237 51
rect -1237 -119 -1203 -85
rect -1237 -187 -1203 -153
rect -1237 -255 -1203 -221
rect -1237 -323 -1203 -289
rect -1237 -391 -1203 -357
rect -1237 -459 -1203 -425
rect -1237 -527 -1203 -493
rect -1237 -595 -1203 -561
rect -1237 -663 -1203 -629
rect -1237 -731 -1203 -697
rect -1237 -799 -1203 -765
rect -1237 -867 -1203 -833
rect -1237 -935 -1203 -901
rect -1237 -1003 -1203 -969
rect -1237 -1071 -1203 -1037
rect -1237 -1139 -1203 -1105
rect -1237 -1207 -1203 -1173
rect -1237 -1275 -1203 -1241
rect 1203 -51 1237 -17
rect 1203 -119 1237 -85
rect 1203 -187 1237 -153
rect 1203 -255 1237 -221
rect 1203 -323 1237 -289
rect 1203 -391 1237 -357
rect 1203 -459 1237 -425
rect 1203 -527 1237 -493
rect 1203 -595 1237 -561
rect 1203 -663 1237 -629
rect 1203 -731 1237 -697
rect 1203 -799 1237 -765
rect 1203 -867 1237 -833
rect 1203 -935 1237 -901
rect 1203 -1003 1237 -969
rect 1203 -1071 1237 -1037
rect 1203 -1139 1237 -1105
rect 1203 -1207 1237 -1173
rect -1237 -1343 -1203 -1309
rect 1203 -1275 1237 -1241
rect 1203 -1343 1237 -1309
rect -1237 -1411 -1203 -1377
rect 1203 -1411 1237 -1377
rect -1237 -1479 -1203 -1445
rect -1237 -1547 -1203 -1513
rect -1237 -1615 -1203 -1581
rect -1237 -1683 -1203 -1649
rect -1237 -1751 -1203 -1717
rect -1237 -1819 -1203 -1785
rect -1237 -1887 -1203 -1853
rect -1237 -1955 -1203 -1921
rect -1237 -2023 -1203 -1989
rect -1237 -2091 -1203 -2057
rect -1237 -2159 -1203 -2125
rect -1237 -2227 -1203 -2193
rect -1237 -2295 -1203 -2261
rect -1237 -2363 -1203 -2329
rect -1237 -2431 -1203 -2397
rect -1237 -2499 -1203 -2465
rect -1237 -2567 -1203 -2533
rect -1237 -2635 -1203 -2601
rect 1203 -1479 1237 -1445
rect 1203 -1547 1237 -1513
rect 1203 -1615 1237 -1581
rect 1203 -1683 1237 -1649
rect 1203 -1751 1237 -1717
rect 1203 -1819 1237 -1785
rect 1203 -1887 1237 -1853
rect 1203 -1955 1237 -1921
rect 1203 -2023 1237 -1989
rect 1203 -2091 1237 -2057
rect 1203 -2159 1237 -2125
rect 1203 -2227 1237 -2193
rect 1203 -2295 1237 -2261
rect 1203 -2363 1237 -2329
rect 1203 -2431 1237 -2397
rect 1203 -2499 1237 -2465
rect 1203 -2567 1237 -2533
rect -1237 -2761 -1203 -2669
rect 1203 -2635 1237 -2601
rect 1203 -2761 1237 -2669
rect -1237 -2795 -1139 -2761
rect -1105 -2795 -1071 -2761
rect -1037 -2795 -1003 -2761
rect -969 -2795 -935 -2761
rect -901 -2795 -867 -2761
rect -833 -2795 -799 -2761
rect -765 -2795 -731 -2761
rect -697 -2795 -663 -2761
rect -629 -2795 -595 -2761
rect -561 -2795 -527 -2761
rect -493 -2795 -459 -2761
rect -425 -2795 -391 -2761
rect -357 -2795 -323 -2761
rect -289 -2795 -255 -2761
rect -221 -2795 -187 -2761
rect -153 -2795 -119 -2761
rect -85 -2795 -51 -2761
rect -17 -2795 17 -2761
rect 51 -2795 85 -2761
rect 119 -2795 153 -2761
rect 187 -2795 221 -2761
rect 255 -2795 289 -2761
rect 323 -2795 357 -2761
rect 391 -2795 425 -2761
rect 459 -2795 493 -2761
rect 527 -2795 561 -2761
rect 595 -2795 629 -2761
rect 663 -2795 697 -2761
rect 731 -2795 765 -2761
rect 799 -2795 833 -2761
rect 867 -2795 901 -2761
rect 935 -2795 969 -2761
rect 1003 -2795 1037 -2761
rect 1071 -2795 1105 -2761
rect 1139 -2795 1237 -2761
<< nsubdiffcont >>
rect -1139 2761 -1105 2795
rect -1071 2761 -1037 2795
rect -1003 2761 -969 2795
rect -935 2761 -901 2795
rect -867 2761 -833 2795
rect -799 2761 -765 2795
rect -731 2761 -697 2795
rect -663 2761 -629 2795
rect -595 2761 -561 2795
rect -527 2761 -493 2795
rect -459 2761 -425 2795
rect -391 2761 -357 2795
rect -323 2761 -289 2795
rect -255 2761 -221 2795
rect -187 2761 -153 2795
rect -119 2761 -85 2795
rect -51 2761 -17 2795
rect 17 2761 51 2795
rect 85 2761 119 2795
rect 153 2761 187 2795
rect 221 2761 255 2795
rect 289 2761 323 2795
rect 357 2761 391 2795
rect 425 2761 459 2795
rect 493 2761 527 2795
rect 561 2761 595 2795
rect 629 2761 663 2795
rect 697 2761 731 2795
rect 765 2761 799 2795
rect 833 2761 867 2795
rect 901 2761 935 2795
rect 969 2761 1003 2795
rect 1037 2761 1071 2795
rect 1105 2761 1139 2795
rect -1237 2635 -1203 2669
rect -1237 2567 -1203 2601
rect -1237 2499 -1203 2533
rect -1237 2431 -1203 2465
rect -1237 2363 -1203 2397
rect -1237 2295 -1203 2329
rect -1237 2227 -1203 2261
rect -1237 2159 -1203 2193
rect -1237 2091 -1203 2125
rect -1237 2023 -1203 2057
rect -1237 1955 -1203 1989
rect -1237 1887 -1203 1921
rect -1237 1819 -1203 1853
rect -1237 1751 -1203 1785
rect -1237 1683 -1203 1717
rect -1237 1615 -1203 1649
rect -1237 1547 -1203 1581
rect -1237 1479 -1203 1513
rect 1203 2635 1237 2669
rect 1203 2567 1237 2601
rect 1203 2499 1237 2533
rect 1203 2431 1237 2465
rect 1203 2363 1237 2397
rect 1203 2295 1237 2329
rect 1203 2227 1237 2261
rect 1203 2159 1237 2193
rect 1203 2091 1237 2125
rect 1203 2023 1237 2057
rect 1203 1955 1237 1989
rect 1203 1887 1237 1921
rect 1203 1819 1237 1853
rect 1203 1751 1237 1785
rect 1203 1683 1237 1717
rect 1203 1615 1237 1649
rect 1203 1547 1237 1581
rect -1237 1411 -1203 1445
rect 1203 1479 1237 1513
rect 1203 1411 1237 1445
rect -1237 1343 -1203 1377
rect 1203 1343 1237 1377
rect -1237 1275 -1203 1309
rect -1237 1207 -1203 1241
rect -1237 1139 -1203 1173
rect -1237 1071 -1203 1105
rect -1237 1003 -1203 1037
rect -1237 935 -1203 969
rect -1237 867 -1203 901
rect -1237 799 -1203 833
rect -1237 731 -1203 765
rect -1237 663 -1203 697
rect -1237 595 -1203 629
rect -1237 527 -1203 561
rect -1237 459 -1203 493
rect -1237 391 -1203 425
rect -1237 323 -1203 357
rect -1237 255 -1203 289
rect -1237 187 -1203 221
rect -1237 119 -1203 153
rect 1203 1275 1237 1309
rect 1203 1207 1237 1241
rect 1203 1139 1237 1173
rect 1203 1071 1237 1105
rect 1203 1003 1237 1037
rect 1203 935 1237 969
rect 1203 867 1237 901
rect 1203 799 1237 833
rect 1203 731 1237 765
rect 1203 663 1237 697
rect 1203 595 1237 629
rect 1203 527 1237 561
rect 1203 459 1237 493
rect 1203 391 1237 425
rect 1203 323 1237 357
rect 1203 255 1237 289
rect 1203 187 1237 221
rect 1203 119 1237 153
rect -1237 51 -1203 85
rect 1203 51 1237 85
rect -1237 -17 -1203 17
rect 1203 -17 1237 17
rect -1237 -85 -1203 -51
rect -1237 -153 -1203 -119
rect -1237 -221 -1203 -187
rect -1237 -289 -1203 -255
rect -1237 -357 -1203 -323
rect -1237 -425 -1203 -391
rect -1237 -493 -1203 -459
rect -1237 -561 -1203 -527
rect -1237 -629 -1203 -595
rect -1237 -697 -1203 -663
rect -1237 -765 -1203 -731
rect -1237 -833 -1203 -799
rect -1237 -901 -1203 -867
rect -1237 -969 -1203 -935
rect -1237 -1037 -1203 -1003
rect -1237 -1105 -1203 -1071
rect -1237 -1173 -1203 -1139
rect -1237 -1241 -1203 -1207
rect 1203 -85 1237 -51
rect 1203 -153 1237 -119
rect 1203 -221 1237 -187
rect 1203 -289 1237 -255
rect 1203 -357 1237 -323
rect 1203 -425 1237 -391
rect 1203 -493 1237 -459
rect 1203 -561 1237 -527
rect 1203 -629 1237 -595
rect 1203 -697 1237 -663
rect 1203 -765 1237 -731
rect 1203 -833 1237 -799
rect 1203 -901 1237 -867
rect 1203 -969 1237 -935
rect 1203 -1037 1237 -1003
rect 1203 -1105 1237 -1071
rect 1203 -1173 1237 -1139
rect 1203 -1241 1237 -1207
rect -1237 -1309 -1203 -1275
rect -1237 -1377 -1203 -1343
rect 1203 -1309 1237 -1275
rect 1203 -1377 1237 -1343
rect -1237 -1445 -1203 -1411
rect -1237 -1513 -1203 -1479
rect -1237 -1581 -1203 -1547
rect -1237 -1649 -1203 -1615
rect -1237 -1717 -1203 -1683
rect -1237 -1785 -1203 -1751
rect -1237 -1853 -1203 -1819
rect -1237 -1921 -1203 -1887
rect -1237 -1989 -1203 -1955
rect -1237 -2057 -1203 -2023
rect -1237 -2125 -1203 -2091
rect -1237 -2193 -1203 -2159
rect -1237 -2261 -1203 -2227
rect -1237 -2329 -1203 -2295
rect -1237 -2397 -1203 -2363
rect -1237 -2465 -1203 -2431
rect -1237 -2533 -1203 -2499
rect -1237 -2601 -1203 -2567
rect 1203 -1445 1237 -1411
rect 1203 -1513 1237 -1479
rect 1203 -1581 1237 -1547
rect 1203 -1649 1237 -1615
rect 1203 -1717 1237 -1683
rect 1203 -1785 1237 -1751
rect 1203 -1853 1237 -1819
rect 1203 -1921 1237 -1887
rect 1203 -1989 1237 -1955
rect 1203 -2057 1237 -2023
rect 1203 -2125 1237 -2091
rect 1203 -2193 1237 -2159
rect 1203 -2261 1237 -2227
rect 1203 -2329 1237 -2295
rect 1203 -2397 1237 -2363
rect 1203 -2465 1237 -2431
rect 1203 -2533 1237 -2499
rect 1203 -2601 1237 -2567
rect -1237 -2669 -1203 -2635
rect 1203 -2669 1237 -2635
rect -1139 -2795 -1105 -2761
rect -1071 -2795 -1037 -2761
rect -1003 -2795 -969 -2761
rect -935 -2795 -901 -2761
rect -867 -2795 -833 -2761
rect -799 -2795 -765 -2761
rect -731 -2795 -697 -2761
rect -663 -2795 -629 -2761
rect -595 -2795 -561 -2761
rect -527 -2795 -493 -2761
rect -459 -2795 -425 -2761
rect -391 -2795 -357 -2761
rect -323 -2795 -289 -2761
rect -255 -2795 -221 -2761
rect -187 -2795 -153 -2761
rect -119 -2795 -85 -2761
rect -51 -2795 -17 -2761
rect 17 -2795 51 -2761
rect 85 -2795 119 -2761
rect 153 -2795 187 -2761
rect 221 -2795 255 -2761
rect 289 -2795 323 -2761
rect 357 -2795 391 -2761
rect 425 -2795 459 -2761
rect 493 -2795 527 -2761
rect 561 -2795 595 -2761
rect 629 -2795 663 -2761
rect 697 -2795 731 -2761
rect 765 -2795 799 -2761
rect 833 -2795 867 -2761
rect 901 -2795 935 -2761
rect 969 -2795 1003 -2761
rect 1037 -2795 1071 -2761
rect 1105 -2795 1139 -2761
<< poly >>
rect -1077 2683 -977 2709
rect -919 2683 -819 2709
rect -761 2683 -661 2709
rect -603 2683 -503 2709
rect -445 2683 -345 2709
rect -287 2683 -187 2709
rect -129 2683 -29 2709
rect 29 2683 129 2709
rect 187 2683 287 2709
rect 345 2683 445 2709
rect 503 2683 603 2709
rect 661 2683 761 2709
rect 819 2683 919 2709
rect 977 2683 1077 2709
rect -1077 1436 -977 1483
rect -1077 1402 -1044 1436
rect -1010 1402 -977 1436
rect -1077 1386 -977 1402
rect -919 1436 -819 1483
rect -919 1402 -886 1436
rect -852 1402 -819 1436
rect -919 1386 -819 1402
rect -761 1436 -661 1483
rect -761 1402 -728 1436
rect -694 1402 -661 1436
rect -761 1386 -661 1402
rect -603 1436 -503 1483
rect -603 1402 -570 1436
rect -536 1402 -503 1436
rect -603 1386 -503 1402
rect -445 1436 -345 1483
rect -445 1402 -412 1436
rect -378 1402 -345 1436
rect -445 1386 -345 1402
rect -287 1436 -187 1483
rect -287 1402 -254 1436
rect -220 1402 -187 1436
rect -287 1386 -187 1402
rect -129 1436 -29 1483
rect -129 1402 -96 1436
rect -62 1402 -29 1436
rect -129 1386 -29 1402
rect 29 1436 129 1483
rect 29 1402 62 1436
rect 96 1402 129 1436
rect 29 1386 129 1402
rect 187 1436 287 1483
rect 187 1402 220 1436
rect 254 1402 287 1436
rect 187 1386 287 1402
rect 345 1436 445 1483
rect 345 1402 378 1436
rect 412 1402 445 1436
rect 345 1386 445 1402
rect 503 1436 603 1483
rect 503 1402 536 1436
rect 570 1402 603 1436
rect 503 1386 603 1402
rect 661 1436 761 1483
rect 661 1402 694 1436
rect 728 1402 761 1436
rect 661 1386 761 1402
rect 819 1436 919 1483
rect 819 1402 852 1436
rect 886 1402 919 1436
rect 819 1386 919 1402
rect 977 1436 1077 1483
rect 977 1402 1010 1436
rect 1044 1402 1077 1436
rect 977 1386 1077 1402
rect -1077 1318 -977 1344
rect -919 1318 -819 1344
rect -761 1318 -661 1344
rect -603 1318 -503 1344
rect -445 1318 -345 1344
rect -287 1318 -187 1344
rect -129 1318 -29 1344
rect 29 1318 129 1344
rect 187 1318 287 1344
rect 345 1318 445 1344
rect 503 1318 603 1344
rect 661 1318 761 1344
rect 819 1318 919 1344
rect 977 1318 1077 1344
rect -1077 71 -977 118
rect -1077 37 -1044 71
rect -1010 37 -977 71
rect -1077 21 -977 37
rect -919 71 -819 118
rect -919 37 -886 71
rect -852 37 -819 71
rect -919 21 -819 37
rect -761 71 -661 118
rect -761 37 -728 71
rect -694 37 -661 71
rect -761 21 -661 37
rect -603 71 -503 118
rect -603 37 -570 71
rect -536 37 -503 71
rect -603 21 -503 37
rect -445 71 -345 118
rect -445 37 -412 71
rect -378 37 -345 71
rect -445 21 -345 37
rect -287 71 -187 118
rect -287 37 -254 71
rect -220 37 -187 71
rect -287 21 -187 37
rect -129 71 -29 118
rect -129 37 -96 71
rect -62 37 -29 71
rect -129 21 -29 37
rect 29 71 129 118
rect 29 37 62 71
rect 96 37 129 71
rect 29 21 129 37
rect 187 71 287 118
rect 187 37 220 71
rect 254 37 287 71
rect 187 21 287 37
rect 345 71 445 118
rect 345 37 378 71
rect 412 37 445 71
rect 345 21 445 37
rect 503 71 603 118
rect 503 37 536 71
rect 570 37 603 71
rect 503 21 603 37
rect 661 71 761 118
rect 661 37 694 71
rect 728 37 761 71
rect 661 21 761 37
rect 819 71 919 118
rect 819 37 852 71
rect 886 37 919 71
rect 819 21 919 37
rect 977 71 1077 118
rect 977 37 1010 71
rect 1044 37 1077 71
rect 977 21 1077 37
rect -1077 -47 -977 -21
rect -919 -47 -819 -21
rect -761 -47 -661 -21
rect -603 -47 -503 -21
rect -445 -47 -345 -21
rect -287 -47 -187 -21
rect -129 -47 -29 -21
rect 29 -47 129 -21
rect 187 -47 287 -21
rect 345 -47 445 -21
rect 503 -47 603 -21
rect 661 -47 761 -21
rect 819 -47 919 -21
rect 977 -47 1077 -21
rect -1077 -1294 -977 -1247
rect -1077 -1328 -1044 -1294
rect -1010 -1328 -977 -1294
rect -1077 -1344 -977 -1328
rect -919 -1294 -819 -1247
rect -919 -1328 -886 -1294
rect -852 -1328 -819 -1294
rect -919 -1344 -819 -1328
rect -761 -1294 -661 -1247
rect -761 -1328 -728 -1294
rect -694 -1328 -661 -1294
rect -761 -1344 -661 -1328
rect -603 -1294 -503 -1247
rect -603 -1328 -570 -1294
rect -536 -1328 -503 -1294
rect -603 -1344 -503 -1328
rect -445 -1294 -345 -1247
rect -445 -1328 -412 -1294
rect -378 -1328 -345 -1294
rect -445 -1344 -345 -1328
rect -287 -1294 -187 -1247
rect -287 -1328 -254 -1294
rect -220 -1328 -187 -1294
rect -287 -1344 -187 -1328
rect -129 -1294 -29 -1247
rect -129 -1328 -96 -1294
rect -62 -1328 -29 -1294
rect -129 -1344 -29 -1328
rect 29 -1294 129 -1247
rect 29 -1328 62 -1294
rect 96 -1328 129 -1294
rect 29 -1344 129 -1328
rect 187 -1294 287 -1247
rect 187 -1328 220 -1294
rect 254 -1328 287 -1294
rect 187 -1344 287 -1328
rect 345 -1294 445 -1247
rect 345 -1328 378 -1294
rect 412 -1328 445 -1294
rect 345 -1344 445 -1328
rect 503 -1294 603 -1247
rect 503 -1328 536 -1294
rect 570 -1328 603 -1294
rect 503 -1344 603 -1328
rect 661 -1294 761 -1247
rect 661 -1328 694 -1294
rect 728 -1328 761 -1294
rect 661 -1344 761 -1328
rect 819 -1294 919 -1247
rect 819 -1328 852 -1294
rect 886 -1328 919 -1294
rect 819 -1344 919 -1328
rect 977 -1294 1077 -1247
rect 977 -1328 1010 -1294
rect 1044 -1328 1077 -1294
rect 977 -1344 1077 -1328
rect -1077 -1412 -977 -1386
rect -919 -1412 -819 -1386
rect -761 -1412 -661 -1386
rect -603 -1412 -503 -1386
rect -445 -1412 -345 -1386
rect -287 -1412 -187 -1386
rect -129 -1412 -29 -1386
rect 29 -1412 129 -1386
rect 187 -1412 287 -1386
rect 345 -1412 445 -1386
rect 503 -1412 603 -1386
rect 661 -1412 761 -1386
rect 819 -1412 919 -1386
rect 977 -1412 1077 -1386
rect -1077 -2659 -977 -2612
rect -1077 -2693 -1044 -2659
rect -1010 -2693 -977 -2659
rect -1077 -2709 -977 -2693
rect -919 -2659 -819 -2612
rect -919 -2693 -886 -2659
rect -852 -2693 -819 -2659
rect -919 -2709 -819 -2693
rect -761 -2659 -661 -2612
rect -761 -2693 -728 -2659
rect -694 -2693 -661 -2659
rect -761 -2709 -661 -2693
rect -603 -2659 -503 -2612
rect -603 -2693 -570 -2659
rect -536 -2693 -503 -2659
rect -603 -2709 -503 -2693
rect -445 -2659 -345 -2612
rect -445 -2693 -412 -2659
rect -378 -2693 -345 -2659
rect -445 -2709 -345 -2693
rect -287 -2659 -187 -2612
rect -287 -2693 -254 -2659
rect -220 -2693 -187 -2659
rect -287 -2709 -187 -2693
rect -129 -2659 -29 -2612
rect -129 -2693 -96 -2659
rect -62 -2693 -29 -2659
rect -129 -2709 -29 -2693
rect 29 -2659 129 -2612
rect 29 -2693 62 -2659
rect 96 -2693 129 -2659
rect 29 -2709 129 -2693
rect 187 -2659 287 -2612
rect 187 -2693 220 -2659
rect 254 -2693 287 -2659
rect 187 -2709 287 -2693
rect 345 -2659 445 -2612
rect 345 -2693 378 -2659
rect 412 -2693 445 -2659
rect 345 -2709 445 -2693
rect 503 -2659 603 -2612
rect 503 -2693 536 -2659
rect 570 -2693 603 -2659
rect 503 -2709 603 -2693
rect 661 -2659 761 -2612
rect 661 -2693 694 -2659
rect 728 -2693 761 -2659
rect 661 -2709 761 -2693
rect 819 -2659 919 -2612
rect 819 -2693 852 -2659
rect 886 -2693 919 -2659
rect 819 -2709 919 -2693
rect 977 -2659 1077 -2612
rect 977 -2693 1010 -2659
rect 1044 -2693 1077 -2659
rect 977 -2709 1077 -2693
<< polycont >>
rect -1044 1402 -1010 1436
rect -886 1402 -852 1436
rect -728 1402 -694 1436
rect -570 1402 -536 1436
rect -412 1402 -378 1436
rect -254 1402 -220 1436
rect -96 1402 -62 1436
rect 62 1402 96 1436
rect 220 1402 254 1436
rect 378 1402 412 1436
rect 536 1402 570 1436
rect 694 1402 728 1436
rect 852 1402 886 1436
rect 1010 1402 1044 1436
rect -1044 37 -1010 71
rect -886 37 -852 71
rect -728 37 -694 71
rect -570 37 -536 71
rect -412 37 -378 71
rect -254 37 -220 71
rect -96 37 -62 71
rect 62 37 96 71
rect 220 37 254 71
rect 378 37 412 71
rect 536 37 570 71
rect 694 37 728 71
rect 852 37 886 71
rect 1010 37 1044 71
rect -1044 -1328 -1010 -1294
rect -886 -1328 -852 -1294
rect -728 -1328 -694 -1294
rect -570 -1328 -536 -1294
rect -412 -1328 -378 -1294
rect -254 -1328 -220 -1294
rect -96 -1328 -62 -1294
rect 62 -1328 96 -1294
rect 220 -1328 254 -1294
rect 378 -1328 412 -1294
rect 536 -1328 570 -1294
rect 694 -1328 728 -1294
rect 852 -1328 886 -1294
rect 1010 -1328 1044 -1294
rect -1044 -2693 -1010 -2659
rect -886 -2693 -852 -2659
rect -728 -2693 -694 -2659
rect -570 -2693 -536 -2659
rect -412 -2693 -378 -2659
rect -254 -2693 -220 -2659
rect -96 -2693 -62 -2659
rect 62 -2693 96 -2659
rect 220 -2693 254 -2659
rect 378 -2693 412 -2659
rect 536 -2693 570 -2659
rect 694 -2693 728 -2659
rect 852 -2693 886 -2659
rect 1010 -2693 1044 -2659
<< locali >>
rect -1237 2761 -1139 2795
rect -1105 2761 -1071 2795
rect -1037 2761 -1003 2795
rect -969 2761 -935 2795
rect -901 2761 -867 2795
rect -833 2761 -799 2795
rect -765 2761 -731 2795
rect -697 2761 -663 2795
rect -629 2761 -595 2795
rect -561 2761 -527 2795
rect -493 2761 -459 2795
rect -425 2761 -391 2795
rect -357 2761 -323 2795
rect -289 2761 -255 2795
rect -221 2761 -187 2795
rect -153 2761 -119 2795
rect -85 2761 -51 2795
rect -17 2761 17 2795
rect 51 2761 85 2795
rect 119 2761 153 2795
rect 187 2761 221 2795
rect 255 2761 289 2795
rect 323 2761 357 2795
rect 391 2761 425 2795
rect 459 2761 493 2795
rect 527 2761 561 2795
rect 595 2761 629 2795
rect 663 2761 697 2795
rect 731 2761 765 2795
rect 799 2761 833 2795
rect 867 2761 901 2795
rect 935 2761 969 2795
rect 1003 2761 1037 2795
rect 1071 2761 1105 2795
rect 1139 2761 1237 2795
rect -1237 2669 -1203 2761
rect -1237 2601 -1203 2635
rect -1237 2533 -1203 2567
rect -1237 2465 -1203 2499
rect -1237 2397 -1203 2431
rect -1237 2329 -1203 2363
rect -1237 2261 -1203 2295
rect -1237 2193 -1203 2227
rect -1237 2125 -1203 2159
rect -1237 2057 -1203 2091
rect -1237 1989 -1203 2023
rect -1237 1921 -1203 1955
rect -1237 1853 -1203 1887
rect -1237 1785 -1203 1819
rect -1237 1717 -1203 1751
rect -1237 1649 -1203 1683
rect -1237 1581 -1203 1615
rect -1237 1513 -1203 1547
rect -1123 2644 -1089 2687
rect -1123 2576 -1089 2606
rect -1123 2508 -1089 2534
rect -1123 2440 -1089 2462
rect -1123 2372 -1089 2390
rect -1123 2304 -1089 2318
rect -1123 2236 -1089 2246
rect -1123 2168 -1089 2174
rect -1123 2100 -1089 2102
rect -1123 2064 -1089 2066
rect -1123 1992 -1089 1998
rect -1123 1920 -1089 1930
rect -1123 1848 -1089 1862
rect -1123 1776 -1089 1794
rect -1123 1704 -1089 1726
rect -1123 1632 -1089 1658
rect -1123 1560 -1089 1590
rect -1123 1479 -1089 1522
rect -965 2644 -931 2687
rect -965 2576 -931 2606
rect -965 2508 -931 2534
rect -965 2440 -931 2462
rect -965 2372 -931 2390
rect -965 2304 -931 2318
rect -965 2236 -931 2246
rect -965 2168 -931 2174
rect -965 2100 -931 2102
rect -965 2064 -931 2066
rect -965 1992 -931 1998
rect -965 1920 -931 1930
rect -965 1848 -931 1862
rect -965 1776 -931 1794
rect -965 1704 -931 1726
rect -965 1632 -931 1658
rect -965 1560 -931 1590
rect -965 1479 -931 1522
rect -807 2644 -773 2687
rect -807 2576 -773 2606
rect -807 2508 -773 2534
rect -807 2440 -773 2462
rect -807 2372 -773 2390
rect -807 2304 -773 2318
rect -807 2236 -773 2246
rect -807 2168 -773 2174
rect -807 2100 -773 2102
rect -807 2064 -773 2066
rect -807 1992 -773 1998
rect -807 1920 -773 1930
rect -807 1848 -773 1862
rect -807 1776 -773 1794
rect -807 1704 -773 1726
rect -807 1632 -773 1658
rect -807 1560 -773 1590
rect -807 1479 -773 1522
rect -649 2644 -615 2687
rect -649 2576 -615 2606
rect -649 2508 -615 2534
rect -649 2440 -615 2462
rect -649 2372 -615 2390
rect -649 2304 -615 2318
rect -649 2236 -615 2246
rect -649 2168 -615 2174
rect -649 2100 -615 2102
rect -649 2064 -615 2066
rect -649 1992 -615 1998
rect -649 1920 -615 1930
rect -649 1848 -615 1862
rect -649 1776 -615 1794
rect -649 1704 -615 1726
rect -649 1632 -615 1658
rect -649 1560 -615 1590
rect -649 1479 -615 1522
rect -491 2644 -457 2687
rect -491 2576 -457 2606
rect -491 2508 -457 2534
rect -491 2440 -457 2462
rect -491 2372 -457 2390
rect -491 2304 -457 2318
rect -491 2236 -457 2246
rect -491 2168 -457 2174
rect -491 2100 -457 2102
rect -491 2064 -457 2066
rect -491 1992 -457 1998
rect -491 1920 -457 1930
rect -491 1848 -457 1862
rect -491 1776 -457 1794
rect -491 1704 -457 1726
rect -491 1632 -457 1658
rect -491 1560 -457 1590
rect -491 1479 -457 1522
rect -333 2644 -299 2687
rect -333 2576 -299 2606
rect -333 2508 -299 2534
rect -333 2440 -299 2462
rect -333 2372 -299 2390
rect -333 2304 -299 2318
rect -333 2236 -299 2246
rect -333 2168 -299 2174
rect -333 2100 -299 2102
rect -333 2064 -299 2066
rect -333 1992 -299 1998
rect -333 1920 -299 1930
rect -333 1848 -299 1862
rect -333 1776 -299 1794
rect -333 1704 -299 1726
rect -333 1632 -299 1658
rect -333 1560 -299 1590
rect -333 1479 -299 1522
rect -175 2644 -141 2687
rect -175 2576 -141 2606
rect -175 2508 -141 2534
rect -175 2440 -141 2462
rect -175 2372 -141 2390
rect -175 2304 -141 2318
rect -175 2236 -141 2246
rect -175 2168 -141 2174
rect -175 2100 -141 2102
rect -175 2064 -141 2066
rect -175 1992 -141 1998
rect -175 1920 -141 1930
rect -175 1848 -141 1862
rect -175 1776 -141 1794
rect -175 1704 -141 1726
rect -175 1632 -141 1658
rect -175 1560 -141 1590
rect -175 1479 -141 1522
rect -17 2644 17 2687
rect -17 2576 17 2606
rect -17 2508 17 2534
rect -17 2440 17 2462
rect -17 2372 17 2390
rect -17 2304 17 2318
rect -17 2236 17 2246
rect -17 2168 17 2174
rect -17 2100 17 2102
rect -17 2064 17 2066
rect -17 1992 17 1998
rect -17 1920 17 1930
rect -17 1848 17 1862
rect -17 1776 17 1794
rect -17 1704 17 1726
rect -17 1632 17 1658
rect -17 1560 17 1590
rect -17 1479 17 1522
rect 141 2644 175 2687
rect 141 2576 175 2606
rect 141 2508 175 2534
rect 141 2440 175 2462
rect 141 2372 175 2390
rect 141 2304 175 2318
rect 141 2236 175 2246
rect 141 2168 175 2174
rect 141 2100 175 2102
rect 141 2064 175 2066
rect 141 1992 175 1998
rect 141 1920 175 1930
rect 141 1848 175 1862
rect 141 1776 175 1794
rect 141 1704 175 1726
rect 141 1632 175 1658
rect 141 1560 175 1590
rect 141 1479 175 1522
rect 299 2644 333 2687
rect 299 2576 333 2606
rect 299 2508 333 2534
rect 299 2440 333 2462
rect 299 2372 333 2390
rect 299 2304 333 2318
rect 299 2236 333 2246
rect 299 2168 333 2174
rect 299 2100 333 2102
rect 299 2064 333 2066
rect 299 1992 333 1998
rect 299 1920 333 1930
rect 299 1848 333 1862
rect 299 1776 333 1794
rect 299 1704 333 1726
rect 299 1632 333 1658
rect 299 1560 333 1590
rect 299 1479 333 1522
rect 457 2644 491 2687
rect 457 2576 491 2606
rect 457 2508 491 2534
rect 457 2440 491 2462
rect 457 2372 491 2390
rect 457 2304 491 2318
rect 457 2236 491 2246
rect 457 2168 491 2174
rect 457 2100 491 2102
rect 457 2064 491 2066
rect 457 1992 491 1998
rect 457 1920 491 1930
rect 457 1848 491 1862
rect 457 1776 491 1794
rect 457 1704 491 1726
rect 457 1632 491 1658
rect 457 1560 491 1590
rect 457 1479 491 1522
rect 615 2644 649 2687
rect 615 2576 649 2606
rect 615 2508 649 2534
rect 615 2440 649 2462
rect 615 2372 649 2390
rect 615 2304 649 2318
rect 615 2236 649 2246
rect 615 2168 649 2174
rect 615 2100 649 2102
rect 615 2064 649 2066
rect 615 1992 649 1998
rect 615 1920 649 1930
rect 615 1848 649 1862
rect 615 1776 649 1794
rect 615 1704 649 1726
rect 615 1632 649 1658
rect 615 1560 649 1590
rect 615 1479 649 1522
rect 773 2644 807 2687
rect 773 2576 807 2606
rect 773 2508 807 2534
rect 773 2440 807 2462
rect 773 2372 807 2390
rect 773 2304 807 2318
rect 773 2236 807 2246
rect 773 2168 807 2174
rect 773 2100 807 2102
rect 773 2064 807 2066
rect 773 1992 807 1998
rect 773 1920 807 1930
rect 773 1848 807 1862
rect 773 1776 807 1794
rect 773 1704 807 1726
rect 773 1632 807 1658
rect 773 1560 807 1590
rect 773 1479 807 1522
rect 931 2644 965 2687
rect 931 2576 965 2606
rect 931 2508 965 2534
rect 931 2440 965 2462
rect 931 2372 965 2390
rect 931 2304 965 2318
rect 931 2236 965 2246
rect 931 2168 965 2174
rect 931 2100 965 2102
rect 931 2064 965 2066
rect 931 1992 965 1998
rect 931 1920 965 1930
rect 931 1848 965 1862
rect 931 1776 965 1794
rect 931 1704 965 1726
rect 931 1632 965 1658
rect 931 1560 965 1590
rect 931 1479 965 1522
rect 1089 2644 1123 2687
rect 1089 2576 1123 2606
rect 1089 2508 1123 2534
rect 1089 2440 1123 2462
rect 1089 2372 1123 2390
rect 1089 2304 1123 2318
rect 1089 2236 1123 2246
rect 1089 2168 1123 2174
rect 1089 2100 1123 2102
rect 1089 2064 1123 2066
rect 1089 1992 1123 1998
rect 1089 1920 1123 1930
rect 1089 1848 1123 1862
rect 1089 1776 1123 1794
rect 1089 1704 1123 1726
rect 1089 1632 1123 1658
rect 1089 1560 1123 1590
rect 1089 1479 1123 1522
rect 1203 2669 1237 2761
rect 1203 2601 1237 2635
rect 1203 2533 1237 2567
rect 1203 2465 1237 2499
rect 1203 2397 1237 2431
rect 1203 2329 1237 2363
rect 1203 2261 1237 2295
rect 1203 2193 1237 2227
rect 1203 2125 1237 2159
rect 1203 2057 1237 2091
rect 1203 1989 1237 2023
rect 1203 1921 1237 1955
rect 1203 1853 1237 1887
rect 1203 1785 1237 1819
rect 1203 1717 1237 1751
rect 1203 1649 1237 1683
rect 1203 1581 1237 1615
rect 1203 1513 1237 1547
rect -1237 1445 -1203 1479
rect 1203 1445 1237 1479
rect -1237 1377 -1203 1411
rect -1077 1402 -1044 1436
rect -1010 1402 -977 1436
rect -919 1402 -886 1436
rect -852 1402 -819 1436
rect -761 1402 -728 1436
rect -694 1402 -661 1436
rect -603 1402 -570 1436
rect -536 1402 -503 1436
rect -445 1402 -412 1436
rect -378 1402 -345 1436
rect -287 1402 -254 1436
rect -220 1402 -187 1436
rect -129 1402 -96 1436
rect -62 1402 -29 1436
rect 29 1402 62 1436
rect 96 1402 129 1436
rect 187 1402 220 1436
rect 254 1402 287 1436
rect 345 1402 378 1436
rect 412 1402 445 1436
rect 503 1402 536 1436
rect 570 1402 603 1436
rect 661 1402 694 1436
rect 728 1402 761 1436
rect 819 1402 852 1436
rect 886 1402 919 1436
rect 977 1402 1010 1436
rect 1044 1402 1077 1436
rect -1237 1309 -1203 1343
rect 1203 1377 1237 1411
rect -1237 1241 -1203 1275
rect -1237 1173 -1203 1207
rect -1237 1105 -1203 1139
rect -1237 1037 -1203 1071
rect -1237 969 -1203 1003
rect -1237 901 -1203 935
rect -1237 833 -1203 867
rect -1237 765 -1203 799
rect -1237 697 -1203 731
rect -1237 629 -1203 663
rect -1237 561 -1203 595
rect -1237 493 -1203 527
rect -1237 425 -1203 459
rect -1237 357 -1203 391
rect -1237 289 -1203 323
rect -1237 221 -1203 255
rect -1237 153 -1203 187
rect -1237 85 -1203 119
rect -1123 1279 -1089 1322
rect -1123 1211 -1089 1241
rect -1123 1143 -1089 1169
rect -1123 1075 -1089 1097
rect -1123 1007 -1089 1025
rect -1123 939 -1089 953
rect -1123 871 -1089 881
rect -1123 803 -1089 809
rect -1123 735 -1089 737
rect -1123 699 -1089 701
rect -1123 627 -1089 633
rect -1123 555 -1089 565
rect -1123 483 -1089 497
rect -1123 411 -1089 429
rect -1123 339 -1089 361
rect -1123 267 -1089 293
rect -1123 195 -1089 225
rect -1123 114 -1089 157
rect -965 1279 -931 1322
rect -965 1211 -931 1241
rect -965 1143 -931 1169
rect -965 1075 -931 1097
rect -965 1007 -931 1025
rect -965 939 -931 953
rect -965 871 -931 881
rect -965 803 -931 809
rect -965 735 -931 737
rect -965 699 -931 701
rect -965 627 -931 633
rect -965 555 -931 565
rect -965 483 -931 497
rect -965 411 -931 429
rect -965 339 -931 361
rect -965 267 -931 293
rect -965 195 -931 225
rect -965 114 -931 157
rect -807 1279 -773 1322
rect -807 1211 -773 1241
rect -807 1143 -773 1169
rect -807 1075 -773 1097
rect -807 1007 -773 1025
rect -807 939 -773 953
rect -807 871 -773 881
rect -807 803 -773 809
rect -807 735 -773 737
rect -807 699 -773 701
rect -807 627 -773 633
rect -807 555 -773 565
rect -807 483 -773 497
rect -807 411 -773 429
rect -807 339 -773 361
rect -807 267 -773 293
rect -807 195 -773 225
rect -807 114 -773 157
rect -649 1279 -615 1322
rect -649 1211 -615 1241
rect -649 1143 -615 1169
rect -649 1075 -615 1097
rect -649 1007 -615 1025
rect -649 939 -615 953
rect -649 871 -615 881
rect -649 803 -615 809
rect -649 735 -615 737
rect -649 699 -615 701
rect -649 627 -615 633
rect -649 555 -615 565
rect -649 483 -615 497
rect -649 411 -615 429
rect -649 339 -615 361
rect -649 267 -615 293
rect -649 195 -615 225
rect -649 114 -615 157
rect -491 1279 -457 1322
rect -491 1211 -457 1241
rect -491 1143 -457 1169
rect -491 1075 -457 1097
rect -491 1007 -457 1025
rect -491 939 -457 953
rect -491 871 -457 881
rect -491 803 -457 809
rect -491 735 -457 737
rect -491 699 -457 701
rect -491 627 -457 633
rect -491 555 -457 565
rect -491 483 -457 497
rect -491 411 -457 429
rect -491 339 -457 361
rect -491 267 -457 293
rect -491 195 -457 225
rect -491 114 -457 157
rect -333 1279 -299 1322
rect -333 1211 -299 1241
rect -333 1143 -299 1169
rect -333 1075 -299 1097
rect -333 1007 -299 1025
rect -333 939 -299 953
rect -333 871 -299 881
rect -333 803 -299 809
rect -333 735 -299 737
rect -333 699 -299 701
rect -333 627 -299 633
rect -333 555 -299 565
rect -333 483 -299 497
rect -333 411 -299 429
rect -333 339 -299 361
rect -333 267 -299 293
rect -333 195 -299 225
rect -333 114 -299 157
rect -175 1279 -141 1322
rect -175 1211 -141 1241
rect -175 1143 -141 1169
rect -175 1075 -141 1097
rect -175 1007 -141 1025
rect -175 939 -141 953
rect -175 871 -141 881
rect -175 803 -141 809
rect -175 735 -141 737
rect -175 699 -141 701
rect -175 627 -141 633
rect -175 555 -141 565
rect -175 483 -141 497
rect -175 411 -141 429
rect -175 339 -141 361
rect -175 267 -141 293
rect -175 195 -141 225
rect -175 114 -141 157
rect -17 1279 17 1322
rect -17 1211 17 1241
rect -17 1143 17 1169
rect -17 1075 17 1097
rect -17 1007 17 1025
rect -17 939 17 953
rect -17 871 17 881
rect -17 803 17 809
rect -17 735 17 737
rect -17 699 17 701
rect -17 627 17 633
rect -17 555 17 565
rect -17 483 17 497
rect -17 411 17 429
rect -17 339 17 361
rect -17 267 17 293
rect -17 195 17 225
rect -17 114 17 157
rect 141 1279 175 1322
rect 141 1211 175 1241
rect 141 1143 175 1169
rect 141 1075 175 1097
rect 141 1007 175 1025
rect 141 939 175 953
rect 141 871 175 881
rect 141 803 175 809
rect 141 735 175 737
rect 141 699 175 701
rect 141 627 175 633
rect 141 555 175 565
rect 141 483 175 497
rect 141 411 175 429
rect 141 339 175 361
rect 141 267 175 293
rect 141 195 175 225
rect 141 114 175 157
rect 299 1279 333 1322
rect 299 1211 333 1241
rect 299 1143 333 1169
rect 299 1075 333 1097
rect 299 1007 333 1025
rect 299 939 333 953
rect 299 871 333 881
rect 299 803 333 809
rect 299 735 333 737
rect 299 699 333 701
rect 299 627 333 633
rect 299 555 333 565
rect 299 483 333 497
rect 299 411 333 429
rect 299 339 333 361
rect 299 267 333 293
rect 299 195 333 225
rect 299 114 333 157
rect 457 1279 491 1322
rect 457 1211 491 1241
rect 457 1143 491 1169
rect 457 1075 491 1097
rect 457 1007 491 1025
rect 457 939 491 953
rect 457 871 491 881
rect 457 803 491 809
rect 457 735 491 737
rect 457 699 491 701
rect 457 627 491 633
rect 457 555 491 565
rect 457 483 491 497
rect 457 411 491 429
rect 457 339 491 361
rect 457 267 491 293
rect 457 195 491 225
rect 457 114 491 157
rect 615 1279 649 1322
rect 615 1211 649 1241
rect 615 1143 649 1169
rect 615 1075 649 1097
rect 615 1007 649 1025
rect 615 939 649 953
rect 615 871 649 881
rect 615 803 649 809
rect 615 735 649 737
rect 615 699 649 701
rect 615 627 649 633
rect 615 555 649 565
rect 615 483 649 497
rect 615 411 649 429
rect 615 339 649 361
rect 615 267 649 293
rect 615 195 649 225
rect 615 114 649 157
rect 773 1279 807 1322
rect 773 1211 807 1241
rect 773 1143 807 1169
rect 773 1075 807 1097
rect 773 1007 807 1025
rect 773 939 807 953
rect 773 871 807 881
rect 773 803 807 809
rect 773 735 807 737
rect 773 699 807 701
rect 773 627 807 633
rect 773 555 807 565
rect 773 483 807 497
rect 773 411 807 429
rect 773 339 807 361
rect 773 267 807 293
rect 773 195 807 225
rect 773 114 807 157
rect 931 1279 965 1322
rect 931 1211 965 1241
rect 931 1143 965 1169
rect 931 1075 965 1097
rect 931 1007 965 1025
rect 931 939 965 953
rect 931 871 965 881
rect 931 803 965 809
rect 931 735 965 737
rect 931 699 965 701
rect 931 627 965 633
rect 931 555 965 565
rect 931 483 965 497
rect 931 411 965 429
rect 931 339 965 361
rect 931 267 965 293
rect 931 195 965 225
rect 931 114 965 157
rect 1089 1279 1123 1322
rect 1089 1211 1123 1241
rect 1089 1143 1123 1169
rect 1089 1075 1123 1097
rect 1089 1007 1123 1025
rect 1089 939 1123 953
rect 1089 871 1123 881
rect 1089 803 1123 809
rect 1089 735 1123 737
rect 1089 699 1123 701
rect 1089 627 1123 633
rect 1089 555 1123 565
rect 1089 483 1123 497
rect 1089 411 1123 429
rect 1089 339 1123 361
rect 1089 267 1123 293
rect 1089 195 1123 225
rect 1089 114 1123 157
rect 1203 1309 1237 1343
rect 1203 1241 1237 1275
rect 1203 1173 1237 1207
rect 1203 1105 1237 1139
rect 1203 1037 1237 1071
rect 1203 969 1237 1003
rect 1203 901 1237 935
rect 1203 833 1237 867
rect 1203 765 1237 799
rect 1203 697 1237 731
rect 1203 629 1237 663
rect 1203 561 1237 595
rect 1203 493 1237 527
rect 1203 425 1237 459
rect 1203 357 1237 391
rect 1203 289 1237 323
rect 1203 221 1237 255
rect 1203 153 1237 187
rect 1203 85 1237 119
rect -1237 17 -1203 51
rect -1077 37 -1044 71
rect -1010 37 -977 71
rect -919 37 -886 71
rect -852 37 -819 71
rect -761 37 -728 71
rect -694 37 -661 71
rect -603 37 -570 71
rect -536 37 -503 71
rect -445 37 -412 71
rect -378 37 -345 71
rect -287 37 -254 71
rect -220 37 -187 71
rect -129 37 -96 71
rect -62 37 -29 71
rect 29 37 62 71
rect 96 37 129 71
rect 187 37 220 71
rect 254 37 287 71
rect 345 37 378 71
rect 412 37 445 71
rect 503 37 536 71
rect 570 37 603 71
rect 661 37 694 71
rect 728 37 761 71
rect 819 37 852 71
rect 886 37 919 71
rect 977 37 1010 71
rect 1044 37 1077 71
rect -1237 -51 -1203 -17
rect 1203 17 1237 51
rect -1237 -119 -1203 -85
rect -1237 -187 -1203 -153
rect -1237 -255 -1203 -221
rect -1237 -323 -1203 -289
rect -1237 -391 -1203 -357
rect -1237 -459 -1203 -425
rect -1237 -527 -1203 -493
rect -1237 -595 -1203 -561
rect -1237 -663 -1203 -629
rect -1237 -731 -1203 -697
rect -1237 -799 -1203 -765
rect -1237 -867 -1203 -833
rect -1237 -935 -1203 -901
rect -1237 -1003 -1203 -969
rect -1237 -1071 -1203 -1037
rect -1237 -1139 -1203 -1105
rect -1237 -1207 -1203 -1173
rect -1237 -1275 -1203 -1241
rect -1123 -86 -1089 -43
rect -1123 -154 -1089 -124
rect -1123 -222 -1089 -196
rect -1123 -290 -1089 -268
rect -1123 -358 -1089 -340
rect -1123 -426 -1089 -412
rect -1123 -494 -1089 -484
rect -1123 -562 -1089 -556
rect -1123 -630 -1089 -628
rect -1123 -666 -1089 -664
rect -1123 -738 -1089 -732
rect -1123 -810 -1089 -800
rect -1123 -882 -1089 -868
rect -1123 -954 -1089 -936
rect -1123 -1026 -1089 -1004
rect -1123 -1098 -1089 -1072
rect -1123 -1170 -1089 -1140
rect -1123 -1251 -1089 -1208
rect -965 -86 -931 -43
rect -965 -154 -931 -124
rect -965 -222 -931 -196
rect -965 -290 -931 -268
rect -965 -358 -931 -340
rect -965 -426 -931 -412
rect -965 -494 -931 -484
rect -965 -562 -931 -556
rect -965 -630 -931 -628
rect -965 -666 -931 -664
rect -965 -738 -931 -732
rect -965 -810 -931 -800
rect -965 -882 -931 -868
rect -965 -954 -931 -936
rect -965 -1026 -931 -1004
rect -965 -1098 -931 -1072
rect -965 -1170 -931 -1140
rect -965 -1251 -931 -1208
rect -807 -86 -773 -43
rect -807 -154 -773 -124
rect -807 -222 -773 -196
rect -807 -290 -773 -268
rect -807 -358 -773 -340
rect -807 -426 -773 -412
rect -807 -494 -773 -484
rect -807 -562 -773 -556
rect -807 -630 -773 -628
rect -807 -666 -773 -664
rect -807 -738 -773 -732
rect -807 -810 -773 -800
rect -807 -882 -773 -868
rect -807 -954 -773 -936
rect -807 -1026 -773 -1004
rect -807 -1098 -773 -1072
rect -807 -1170 -773 -1140
rect -807 -1251 -773 -1208
rect -649 -86 -615 -43
rect -649 -154 -615 -124
rect -649 -222 -615 -196
rect -649 -290 -615 -268
rect -649 -358 -615 -340
rect -649 -426 -615 -412
rect -649 -494 -615 -484
rect -649 -562 -615 -556
rect -649 -630 -615 -628
rect -649 -666 -615 -664
rect -649 -738 -615 -732
rect -649 -810 -615 -800
rect -649 -882 -615 -868
rect -649 -954 -615 -936
rect -649 -1026 -615 -1004
rect -649 -1098 -615 -1072
rect -649 -1170 -615 -1140
rect -649 -1251 -615 -1208
rect -491 -86 -457 -43
rect -491 -154 -457 -124
rect -491 -222 -457 -196
rect -491 -290 -457 -268
rect -491 -358 -457 -340
rect -491 -426 -457 -412
rect -491 -494 -457 -484
rect -491 -562 -457 -556
rect -491 -630 -457 -628
rect -491 -666 -457 -664
rect -491 -738 -457 -732
rect -491 -810 -457 -800
rect -491 -882 -457 -868
rect -491 -954 -457 -936
rect -491 -1026 -457 -1004
rect -491 -1098 -457 -1072
rect -491 -1170 -457 -1140
rect -491 -1251 -457 -1208
rect -333 -86 -299 -43
rect -333 -154 -299 -124
rect -333 -222 -299 -196
rect -333 -290 -299 -268
rect -333 -358 -299 -340
rect -333 -426 -299 -412
rect -333 -494 -299 -484
rect -333 -562 -299 -556
rect -333 -630 -299 -628
rect -333 -666 -299 -664
rect -333 -738 -299 -732
rect -333 -810 -299 -800
rect -333 -882 -299 -868
rect -333 -954 -299 -936
rect -333 -1026 -299 -1004
rect -333 -1098 -299 -1072
rect -333 -1170 -299 -1140
rect -333 -1251 -299 -1208
rect -175 -86 -141 -43
rect -175 -154 -141 -124
rect -175 -222 -141 -196
rect -175 -290 -141 -268
rect -175 -358 -141 -340
rect -175 -426 -141 -412
rect -175 -494 -141 -484
rect -175 -562 -141 -556
rect -175 -630 -141 -628
rect -175 -666 -141 -664
rect -175 -738 -141 -732
rect -175 -810 -141 -800
rect -175 -882 -141 -868
rect -175 -954 -141 -936
rect -175 -1026 -141 -1004
rect -175 -1098 -141 -1072
rect -175 -1170 -141 -1140
rect -175 -1251 -141 -1208
rect -17 -86 17 -43
rect -17 -154 17 -124
rect -17 -222 17 -196
rect -17 -290 17 -268
rect -17 -358 17 -340
rect -17 -426 17 -412
rect -17 -494 17 -484
rect -17 -562 17 -556
rect -17 -630 17 -628
rect -17 -666 17 -664
rect -17 -738 17 -732
rect -17 -810 17 -800
rect -17 -882 17 -868
rect -17 -954 17 -936
rect -17 -1026 17 -1004
rect -17 -1098 17 -1072
rect -17 -1170 17 -1140
rect -17 -1251 17 -1208
rect 141 -86 175 -43
rect 141 -154 175 -124
rect 141 -222 175 -196
rect 141 -290 175 -268
rect 141 -358 175 -340
rect 141 -426 175 -412
rect 141 -494 175 -484
rect 141 -562 175 -556
rect 141 -630 175 -628
rect 141 -666 175 -664
rect 141 -738 175 -732
rect 141 -810 175 -800
rect 141 -882 175 -868
rect 141 -954 175 -936
rect 141 -1026 175 -1004
rect 141 -1098 175 -1072
rect 141 -1170 175 -1140
rect 141 -1251 175 -1208
rect 299 -86 333 -43
rect 299 -154 333 -124
rect 299 -222 333 -196
rect 299 -290 333 -268
rect 299 -358 333 -340
rect 299 -426 333 -412
rect 299 -494 333 -484
rect 299 -562 333 -556
rect 299 -630 333 -628
rect 299 -666 333 -664
rect 299 -738 333 -732
rect 299 -810 333 -800
rect 299 -882 333 -868
rect 299 -954 333 -936
rect 299 -1026 333 -1004
rect 299 -1098 333 -1072
rect 299 -1170 333 -1140
rect 299 -1251 333 -1208
rect 457 -86 491 -43
rect 457 -154 491 -124
rect 457 -222 491 -196
rect 457 -290 491 -268
rect 457 -358 491 -340
rect 457 -426 491 -412
rect 457 -494 491 -484
rect 457 -562 491 -556
rect 457 -630 491 -628
rect 457 -666 491 -664
rect 457 -738 491 -732
rect 457 -810 491 -800
rect 457 -882 491 -868
rect 457 -954 491 -936
rect 457 -1026 491 -1004
rect 457 -1098 491 -1072
rect 457 -1170 491 -1140
rect 457 -1251 491 -1208
rect 615 -86 649 -43
rect 615 -154 649 -124
rect 615 -222 649 -196
rect 615 -290 649 -268
rect 615 -358 649 -340
rect 615 -426 649 -412
rect 615 -494 649 -484
rect 615 -562 649 -556
rect 615 -630 649 -628
rect 615 -666 649 -664
rect 615 -738 649 -732
rect 615 -810 649 -800
rect 615 -882 649 -868
rect 615 -954 649 -936
rect 615 -1026 649 -1004
rect 615 -1098 649 -1072
rect 615 -1170 649 -1140
rect 615 -1251 649 -1208
rect 773 -86 807 -43
rect 773 -154 807 -124
rect 773 -222 807 -196
rect 773 -290 807 -268
rect 773 -358 807 -340
rect 773 -426 807 -412
rect 773 -494 807 -484
rect 773 -562 807 -556
rect 773 -630 807 -628
rect 773 -666 807 -664
rect 773 -738 807 -732
rect 773 -810 807 -800
rect 773 -882 807 -868
rect 773 -954 807 -936
rect 773 -1026 807 -1004
rect 773 -1098 807 -1072
rect 773 -1170 807 -1140
rect 773 -1251 807 -1208
rect 931 -86 965 -43
rect 931 -154 965 -124
rect 931 -222 965 -196
rect 931 -290 965 -268
rect 931 -358 965 -340
rect 931 -426 965 -412
rect 931 -494 965 -484
rect 931 -562 965 -556
rect 931 -630 965 -628
rect 931 -666 965 -664
rect 931 -738 965 -732
rect 931 -810 965 -800
rect 931 -882 965 -868
rect 931 -954 965 -936
rect 931 -1026 965 -1004
rect 931 -1098 965 -1072
rect 931 -1170 965 -1140
rect 931 -1251 965 -1208
rect 1089 -86 1123 -43
rect 1089 -154 1123 -124
rect 1089 -222 1123 -196
rect 1089 -290 1123 -268
rect 1089 -358 1123 -340
rect 1089 -426 1123 -412
rect 1089 -494 1123 -484
rect 1089 -562 1123 -556
rect 1089 -630 1123 -628
rect 1089 -666 1123 -664
rect 1089 -738 1123 -732
rect 1089 -810 1123 -800
rect 1089 -882 1123 -868
rect 1089 -954 1123 -936
rect 1089 -1026 1123 -1004
rect 1089 -1098 1123 -1072
rect 1089 -1170 1123 -1140
rect 1089 -1251 1123 -1208
rect 1203 -51 1237 -17
rect 1203 -119 1237 -85
rect 1203 -187 1237 -153
rect 1203 -255 1237 -221
rect 1203 -323 1237 -289
rect 1203 -391 1237 -357
rect 1203 -459 1237 -425
rect 1203 -527 1237 -493
rect 1203 -595 1237 -561
rect 1203 -663 1237 -629
rect 1203 -731 1237 -697
rect 1203 -799 1237 -765
rect 1203 -867 1237 -833
rect 1203 -935 1237 -901
rect 1203 -1003 1237 -969
rect 1203 -1071 1237 -1037
rect 1203 -1139 1237 -1105
rect 1203 -1207 1237 -1173
rect 1203 -1275 1237 -1241
rect -1237 -1343 -1203 -1309
rect -1077 -1328 -1044 -1294
rect -1010 -1328 -977 -1294
rect -919 -1328 -886 -1294
rect -852 -1328 -819 -1294
rect -761 -1328 -728 -1294
rect -694 -1328 -661 -1294
rect -603 -1328 -570 -1294
rect -536 -1328 -503 -1294
rect -445 -1328 -412 -1294
rect -378 -1328 -345 -1294
rect -287 -1328 -254 -1294
rect -220 -1328 -187 -1294
rect -129 -1328 -96 -1294
rect -62 -1328 -29 -1294
rect 29 -1328 62 -1294
rect 96 -1328 129 -1294
rect 187 -1328 220 -1294
rect 254 -1328 287 -1294
rect 345 -1328 378 -1294
rect 412 -1328 445 -1294
rect 503 -1328 536 -1294
rect 570 -1328 603 -1294
rect 661 -1328 694 -1294
rect 728 -1328 761 -1294
rect 819 -1328 852 -1294
rect 886 -1328 919 -1294
rect 977 -1328 1010 -1294
rect 1044 -1328 1077 -1294
rect -1237 -1411 -1203 -1377
rect 1203 -1343 1237 -1309
rect -1237 -1479 -1203 -1445
rect -1237 -1547 -1203 -1513
rect -1237 -1615 -1203 -1581
rect -1237 -1683 -1203 -1649
rect -1237 -1751 -1203 -1717
rect -1237 -1819 -1203 -1785
rect -1237 -1887 -1203 -1853
rect -1237 -1955 -1203 -1921
rect -1237 -2023 -1203 -1989
rect -1237 -2091 -1203 -2057
rect -1237 -2159 -1203 -2125
rect -1237 -2227 -1203 -2193
rect -1237 -2295 -1203 -2261
rect -1237 -2363 -1203 -2329
rect -1237 -2431 -1203 -2397
rect -1237 -2499 -1203 -2465
rect -1237 -2567 -1203 -2533
rect -1237 -2635 -1203 -2601
rect -1123 -1451 -1089 -1408
rect -1123 -1519 -1089 -1489
rect -1123 -1587 -1089 -1561
rect -1123 -1655 -1089 -1633
rect -1123 -1723 -1089 -1705
rect -1123 -1791 -1089 -1777
rect -1123 -1859 -1089 -1849
rect -1123 -1927 -1089 -1921
rect -1123 -1995 -1089 -1993
rect -1123 -2031 -1089 -2029
rect -1123 -2103 -1089 -2097
rect -1123 -2175 -1089 -2165
rect -1123 -2247 -1089 -2233
rect -1123 -2319 -1089 -2301
rect -1123 -2391 -1089 -2369
rect -1123 -2463 -1089 -2437
rect -1123 -2535 -1089 -2505
rect -1123 -2616 -1089 -2573
rect -965 -1451 -931 -1408
rect -965 -1519 -931 -1489
rect -965 -1587 -931 -1561
rect -965 -1655 -931 -1633
rect -965 -1723 -931 -1705
rect -965 -1791 -931 -1777
rect -965 -1859 -931 -1849
rect -965 -1927 -931 -1921
rect -965 -1995 -931 -1993
rect -965 -2031 -931 -2029
rect -965 -2103 -931 -2097
rect -965 -2175 -931 -2165
rect -965 -2247 -931 -2233
rect -965 -2319 -931 -2301
rect -965 -2391 -931 -2369
rect -965 -2463 -931 -2437
rect -965 -2535 -931 -2505
rect -965 -2616 -931 -2573
rect -807 -1451 -773 -1408
rect -807 -1519 -773 -1489
rect -807 -1587 -773 -1561
rect -807 -1655 -773 -1633
rect -807 -1723 -773 -1705
rect -807 -1791 -773 -1777
rect -807 -1859 -773 -1849
rect -807 -1927 -773 -1921
rect -807 -1995 -773 -1993
rect -807 -2031 -773 -2029
rect -807 -2103 -773 -2097
rect -807 -2175 -773 -2165
rect -807 -2247 -773 -2233
rect -807 -2319 -773 -2301
rect -807 -2391 -773 -2369
rect -807 -2463 -773 -2437
rect -807 -2535 -773 -2505
rect -807 -2616 -773 -2573
rect -649 -1451 -615 -1408
rect -649 -1519 -615 -1489
rect -649 -1587 -615 -1561
rect -649 -1655 -615 -1633
rect -649 -1723 -615 -1705
rect -649 -1791 -615 -1777
rect -649 -1859 -615 -1849
rect -649 -1927 -615 -1921
rect -649 -1995 -615 -1993
rect -649 -2031 -615 -2029
rect -649 -2103 -615 -2097
rect -649 -2175 -615 -2165
rect -649 -2247 -615 -2233
rect -649 -2319 -615 -2301
rect -649 -2391 -615 -2369
rect -649 -2463 -615 -2437
rect -649 -2535 -615 -2505
rect -649 -2616 -615 -2573
rect -491 -1451 -457 -1408
rect -491 -1519 -457 -1489
rect -491 -1587 -457 -1561
rect -491 -1655 -457 -1633
rect -491 -1723 -457 -1705
rect -491 -1791 -457 -1777
rect -491 -1859 -457 -1849
rect -491 -1927 -457 -1921
rect -491 -1995 -457 -1993
rect -491 -2031 -457 -2029
rect -491 -2103 -457 -2097
rect -491 -2175 -457 -2165
rect -491 -2247 -457 -2233
rect -491 -2319 -457 -2301
rect -491 -2391 -457 -2369
rect -491 -2463 -457 -2437
rect -491 -2535 -457 -2505
rect -491 -2616 -457 -2573
rect -333 -1451 -299 -1408
rect -333 -1519 -299 -1489
rect -333 -1587 -299 -1561
rect -333 -1655 -299 -1633
rect -333 -1723 -299 -1705
rect -333 -1791 -299 -1777
rect -333 -1859 -299 -1849
rect -333 -1927 -299 -1921
rect -333 -1995 -299 -1993
rect -333 -2031 -299 -2029
rect -333 -2103 -299 -2097
rect -333 -2175 -299 -2165
rect -333 -2247 -299 -2233
rect -333 -2319 -299 -2301
rect -333 -2391 -299 -2369
rect -333 -2463 -299 -2437
rect -333 -2535 -299 -2505
rect -333 -2616 -299 -2573
rect -175 -1451 -141 -1408
rect -175 -1519 -141 -1489
rect -175 -1587 -141 -1561
rect -175 -1655 -141 -1633
rect -175 -1723 -141 -1705
rect -175 -1791 -141 -1777
rect -175 -1859 -141 -1849
rect -175 -1927 -141 -1921
rect -175 -1995 -141 -1993
rect -175 -2031 -141 -2029
rect -175 -2103 -141 -2097
rect -175 -2175 -141 -2165
rect -175 -2247 -141 -2233
rect -175 -2319 -141 -2301
rect -175 -2391 -141 -2369
rect -175 -2463 -141 -2437
rect -175 -2535 -141 -2505
rect -175 -2616 -141 -2573
rect -17 -1451 17 -1408
rect -17 -1519 17 -1489
rect -17 -1587 17 -1561
rect -17 -1655 17 -1633
rect -17 -1723 17 -1705
rect -17 -1791 17 -1777
rect -17 -1859 17 -1849
rect -17 -1927 17 -1921
rect -17 -1995 17 -1993
rect -17 -2031 17 -2029
rect -17 -2103 17 -2097
rect -17 -2175 17 -2165
rect -17 -2247 17 -2233
rect -17 -2319 17 -2301
rect -17 -2391 17 -2369
rect -17 -2463 17 -2437
rect -17 -2535 17 -2505
rect -17 -2616 17 -2573
rect 141 -1451 175 -1408
rect 141 -1519 175 -1489
rect 141 -1587 175 -1561
rect 141 -1655 175 -1633
rect 141 -1723 175 -1705
rect 141 -1791 175 -1777
rect 141 -1859 175 -1849
rect 141 -1927 175 -1921
rect 141 -1995 175 -1993
rect 141 -2031 175 -2029
rect 141 -2103 175 -2097
rect 141 -2175 175 -2165
rect 141 -2247 175 -2233
rect 141 -2319 175 -2301
rect 141 -2391 175 -2369
rect 141 -2463 175 -2437
rect 141 -2535 175 -2505
rect 141 -2616 175 -2573
rect 299 -1451 333 -1408
rect 299 -1519 333 -1489
rect 299 -1587 333 -1561
rect 299 -1655 333 -1633
rect 299 -1723 333 -1705
rect 299 -1791 333 -1777
rect 299 -1859 333 -1849
rect 299 -1927 333 -1921
rect 299 -1995 333 -1993
rect 299 -2031 333 -2029
rect 299 -2103 333 -2097
rect 299 -2175 333 -2165
rect 299 -2247 333 -2233
rect 299 -2319 333 -2301
rect 299 -2391 333 -2369
rect 299 -2463 333 -2437
rect 299 -2535 333 -2505
rect 299 -2616 333 -2573
rect 457 -1451 491 -1408
rect 457 -1519 491 -1489
rect 457 -1587 491 -1561
rect 457 -1655 491 -1633
rect 457 -1723 491 -1705
rect 457 -1791 491 -1777
rect 457 -1859 491 -1849
rect 457 -1927 491 -1921
rect 457 -1995 491 -1993
rect 457 -2031 491 -2029
rect 457 -2103 491 -2097
rect 457 -2175 491 -2165
rect 457 -2247 491 -2233
rect 457 -2319 491 -2301
rect 457 -2391 491 -2369
rect 457 -2463 491 -2437
rect 457 -2535 491 -2505
rect 457 -2616 491 -2573
rect 615 -1451 649 -1408
rect 615 -1519 649 -1489
rect 615 -1587 649 -1561
rect 615 -1655 649 -1633
rect 615 -1723 649 -1705
rect 615 -1791 649 -1777
rect 615 -1859 649 -1849
rect 615 -1927 649 -1921
rect 615 -1995 649 -1993
rect 615 -2031 649 -2029
rect 615 -2103 649 -2097
rect 615 -2175 649 -2165
rect 615 -2247 649 -2233
rect 615 -2319 649 -2301
rect 615 -2391 649 -2369
rect 615 -2463 649 -2437
rect 615 -2535 649 -2505
rect 615 -2616 649 -2573
rect 773 -1451 807 -1408
rect 773 -1519 807 -1489
rect 773 -1587 807 -1561
rect 773 -1655 807 -1633
rect 773 -1723 807 -1705
rect 773 -1791 807 -1777
rect 773 -1859 807 -1849
rect 773 -1927 807 -1921
rect 773 -1995 807 -1993
rect 773 -2031 807 -2029
rect 773 -2103 807 -2097
rect 773 -2175 807 -2165
rect 773 -2247 807 -2233
rect 773 -2319 807 -2301
rect 773 -2391 807 -2369
rect 773 -2463 807 -2437
rect 773 -2535 807 -2505
rect 773 -2616 807 -2573
rect 931 -1451 965 -1408
rect 931 -1519 965 -1489
rect 931 -1587 965 -1561
rect 931 -1655 965 -1633
rect 931 -1723 965 -1705
rect 931 -1791 965 -1777
rect 931 -1859 965 -1849
rect 931 -1927 965 -1921
rect 931 -1995 965 -1993
rect 931 -2031 965 -2029
rect 931 -2103 965 -2097
rect 931 -2175 965 -2165
rect 931 -2247 965 -2233
rect 931 -2319 965 -2301
rect 931 -2391 965 -2369
rect 931 -2463 965 -2437
rect 931 -2535 965 -2505
rect 931 -2616 965 -2573
rect 1089 -1451 1123 -1408
rect 1089 -1519 1123 -1489
rect 1089 -1587 1123 -1561
rect 1089 -1655 1123 -1633
rect 1089 -1723 1123 -1705
rect 1089 -1791 1123 -1777
rect 1089 -1859 1123 -1849
rect 1089 -1927 1123 -1921
rect 1089 -1995 1123 -1993
rect 1089 -2031 1123 -2029
rect 1089 -2103 1123 -2097
rect 1089 -2175 1123 -2165
rect 1089 -2247 1123 -2233
rect 1089 -2319 1123 -2301
rect 1089 -2391 1123 -2369
rect 1089 -2463 1123 -2437
rect 1089 -2535 1123 -2505
rect 1089 -2616 1123 -2573
rect 1203 -1411 1237 -1377
rect 1203 -1479 1237 -1445
rect 1203 -1547 1237 -1513
rect 1203 -1615 1237 -1581
rect 1203 -1683 1237 -1649
rect 1203 -1751 1237 -1717
rect 1203 -1819 1237 -1785
rect 1203 -1887 1237 -1853
rect 1203 -1955 1237 -1921
rect 1203 -2023 1237 -1989
rect 1203 -2091 1237 -2057
rect 1203 -2159 1237 -2125
rect 1203 -2227 1237 -2193
rect 1203 -2295 1237 -2261
rect 1203 -2363 1237 -2329
rect 1203 -2431 1237 -2397
rect 1203 -2499 1237 -2465
rect 1203 -2567 1237 -2533
rect 1203 -2635 1237 -2601
rect -1237 -2761 -1203 -2669
rect -1077 -2693 -1044 -2659
rect -1010 -2693 -977 -2659
rect -919 -2693 -886 -2659
rect -852 -2693 -819 -2659
rect -761 -2693 -728 -2659
rect -694 -2693 -661 -2659
rect -603 -2693 -570 -2659
rect -536 -2693 -503 -2659
rect -445 -2693 -412 -2659
rect -378 -2693 -345 -2659
rect -287 -2693 -254 -2659
rect -220 -2693 -187 -2659
rect -129 -2693 -96 -2659
rect -62 -2693 -29 -2659
rect 29 -2693 62 -2659
rect 96 -2693 129 -2659
rect 187 -2693 220 -2659
rect 254 -2693 287 -2659
rect 345 -2693 378 -2659
rect 412 -2693 445 -2659
rect 503 -2693 536 -2659
rect 570 -2693 603 -2659
rect 661 -2693 694 -2659
rect 728 -2693 761 -2659
rect 819 -2693 852 -2659
rect 886 -2693 919 -2659
rect 977 -2693 1010 -2659
rect 1044 -2693 1077 -2659
rect 1203 -2761 1237 -2669
rect -1237 -2795 -1139 -2761
rect -1105 -2795 -1071 -2761
rect -1037 -2795 -1003 -2761
rect -969 -2795 -935 -2761
rect -901 -2795 -867 -2761
rect -833 -2795 -799 -2761
rect -765 -2795 -731 -2761
rect -697 -2795 -663 -2761
rect -629 -2795 -595 -2761
rect -561 -2795 -527 -2761
rect -493 -2795 -459 -2761
rect -425 -2795 -391 -2761
rect -357 -2795 -323 -2761
rect -289 -2795 -255 -2761
rect -221 -2795 -187 -2761
rect -153 -2795 -119 -2761
rect -85 -2795 -51 -2761
rect -17 -2795 17 -2761
rect 51 -2795 85 -2761
rect 119 -2795 153 -2761
rect 187 -2795 221 -2761
rect 255 -2795 289 -2761
rect 323 -2795 357 -2761
rect 391 -2795 425 -2761
rect 459 -2795 493 -2761
rect 527 -2795 561 -2761
rect 595 -2795 629 -2761
rect 663 -2795 697 -2761
rect 731 -2795 765 -2761
rect 799 -2795 833 -2761
rect 867 -2795 901 -2761
rect 935 -2795 969 -2761
rect 1003 -2795 1037 -2761
rect 1071 -2795 1105 -2761
rect 1139 -2795 1237 -2761
<< viali >>
rect -1123 2610 -1089 2640
rect -1123 2606 -1089 2610
rect -1123 2542 -1089 2568
rect -1123 2534 -1089 2542
rect -1123 2474 -1089 2496
rect -1123 2462 -1089 2474
rect -1123 2406 -1089 2424
rect -1123 2390 -1089 2406
rect -1123 2338 -1089 2352
rect -1123 2318 -1089 2338
rect -1123 2270 -1089 2280
rect -1123 2246 -1089 2270
rect -1123 2202 -1089 2208
rect -1123 2174 -1089 2202
rect -1123 2134 -1089 2136
rect -1123 2102 -1089 2134
rect -1123 2032 -1089 2064
rect -1123 2030 -1089 2032
rect -1123 1964 -1089 1992
rect -1123 1958 -1089 1964
rect -1123 1896 -1089 1920
rect -1123 1886 -1089 1896
rect -1123 1828 -1089 1848
rect -1123 1814 -1089 1828
rect -1123 1760 -1089 1776
rect -1123 1742 -1089 1760
rect -1123 1692 -1089 1704
rect -1123 1670 -1089 1692
rect -1123 1624 -1089 1632
rect -1123 1598 -1089 1624
rect -1123 1556 -1089 1560
rect -1123 1526 -1089 1556
rect -965 2610 -931 2640
rect -965 2606 -931 2610
rect -965 2542 -931 2568
rect -965 2534 -931 2542
rect -965 2474 -931 2496
rect -965 2462 -931 2474
rect -965 2406 -931 2424
rect -965 2390 -931 2406
rect -965 2338 -931 2352
rect -965 2318 -931 2338
rect -965 2270 -931 2280
rect -965 2246 -931 2270
rect -965 2202 -931 2208
rect -965 2174 -931 2202
rect -965 2134 -931 2136
rect -965 2102 -931 2134
rect -965 2032 -931 2064
rect -965 2030 -931 2032
rect -965 1964 -931 1992
rect -965 1958 -931 1964
rect -965 1896 -931 1920
rect -965 1886 -931 1896
rect -965 1828 -931 1848
rect -965 1814 -931 1828
rect -965 1760 -931 1776
rect -965 1742 -931 1760
rect -965 1692 -931 1704
rect -965 1670 -931 1692
rect -965 1624 -931 1632
rect -965 1598 -931 1624
rect -965 1556 -931 1560
rect -965 1526 -931 1556
rect -807 2610 -773 2640
rect -807 2606 -773 2610
rect -807 2542 -773 2568
rect -807 2534 -773 2542
rect -807 2474 -773 2496
rect -807 2462 -773 2474
rect -807 2406 -773 2424
rect -807 2390 -773 2406
rect -807 2338 -773 2352
rect -807 2318 -773 2338
rect -807 2270 -773 2280
rect -807 2246 -773 2270
rect -807 2202 -773 2208
rect -807 2174 -773 2202
rect -807 2134 -773 2136
rect -807 2102 -773 2134
rect -807 2032 -773 2064
rect -807 2030 -773 2032
rect -807 1964 -773 1992
rect -807 1958 -773 1964
rect -807 1896 -773 1920
rect -807 1886 -773 1896
rect -807 1828 -773 1848
rect -807 1814 -773 1828
rect -807 1760 -773 1776
rect -807 1742 -773 1760
rect -807 1692 -773 1704
rect -807 1670 -773 1692
rect -807 1624 -773 1632
rect -807 1598 -773 1624
rect -807 1556 -773 1560
rect -807 1526 -773 1556
rect -649 2610 -615 2640
rect -649 2606 -615 2610
rect -649 2542 -615 2568
rect -649 2534 -615 2542
rect -649 2474 -615 2496
rect -649 2462 -615 2474
rect -649 2406 -615 2424
rect -649 2390 -615 2406
rect -649 2338 -615 2352
rect -649 2318 -615 2338
rect -649 2270 -615 2280
rect -649 2246 -615 2270
rect -649 2202 -615 2208
rect -649 2174 -615 2202
rect -649 2134 -615 2136
rect -649 2102 -615 2134
rect -649 2032 -615 2064
rect -649 2030 -615 2032
rect -649 1964 -615 1992
rect -649 1958 -615 1964
rect -649 1896 -615 1920
rect -649 1886 -615 1896
rect -649 1828 -615 1848
rect -649 1814 -615 1828
rect -649 1760 -615 1776
rect -649 1742 -615 1760
rect -649 1692 -615 1704
rect -649 1670 -615 1692
rect -649 1624 -615 1632
rect -649 1598 -615 1624
rect -649 1556 -615 1560
rect -649 1526 -615 1556
rect -491 2610 -457 2640
rect -491 2606 -457 2610
rect -491 2542 -457 2568
rect -491 2534 -457 2542
rect -491 2474 -457 2496
rect -491 2462 -457 2474
rect -491 2406 -457 2424
rect -491 2390 -457 2406
rect -491 2338 -457 2352
rect -491 2318 -457 2338
rect -491 2270 -457 2280
rect -491 2246 -457 2270
rect -491 2202 -457 2208
rect -491 2174 -457 2202
rect -491 2134 -457 2136
rect -491 2102 -457 2134
rect -491 2032 -457 2064
rect -491 2030 -457 2032
rect -491 1964 -457 1992
rect -491 1958 -457 1964
rect -491 1896 -457 1920
rect -491 1886 -457 1896
rect -491 1828 -457 1848
rect -491 1814 -457 1828
rect -491 1760 -457 1776
rect -491 1742 -457 1760
rect -491 1692 -457 1704
rect -491 1670 -457 1692
rect -491 1624 -457 1632
rect -491 1598 -457 1624
rect -491 1556 -457 1560
rect -491 1526 -457 1556
rect -333 2610 -299 2640
rect -333 2606 -299 2610
rect -333 2542 -299 2568
rect -333 2534 -299 2542
rect -333 2474 -299 2496
rect -333 2462 -299 2474
rect -333 2406 -299 2424
rect -333 2390 -299 2406
rect -333 2338 -299 2352
rect -333 2318 -299 2338
rect -333 2270 -299 2280
rect -333 2246 -299 2270
rect -333 2202 -299 2208
rect -333 2174 -299 2202
rect -333 2134 -299 2136
rect -333 2102 -299 2134
rect -333 2032 -299 2064
rect -333 2030 -299 2032
rect -333 1964 -299 1992
rect -333 1958 -299 1964
rect -333 1896 -299 1920
rect -333 1886 -299 1896
rect -333 1828 -299 1848
rect -333 1814 -299 1828
rect -333 1760 -299 1776
rect -333 1742 -299 1760
rect -333 1692 -299 1704
rect -333 1670 -299 1692
rect -333 1624 -299 1632
rect -333 1598 -299 1624
rect -333 1556 -299 1560
rect -333 1526 -299 1556
rect -175 2610 -141 2640
rect -175 2606 -141 2610
rect -175 2542 -141 2568
rect -175 2534 -141 2542
rect -175 2474 -141 2496
rect -175 2462 -141 2474
rect -175 2406 -141 2424
rect -175 2390 -141 2406
rect -175 2338 -141 2352
rect -175 2318 -141 2338
rect -175 2270 -141 2280
rect -175 2246 -141 2270
rect -175 2202 -141 2208
rect -175 2174 -141 2202
rect -175 2134 -141 2136
rect -175 2102 -141 2134
rect -175 2032 -141 2064
rect -175 2030 -141 2032
rect -175 1964 -141 1992
rect -175 1958 -141 1964
rect -175 1896 -141 1920
rect -175 1886 -141 1896
rect -175 1828 -141 1848
rect -175 1814 -141 1828
rect -175 1760 -141 1776
rect -175 1742 -141 1760
rect -175 1692 -141 1704
rect -175 1670 -141 1692
rect -175 1624 -141 1632
rect -175 1598 -141 1624
rect -175 1556 -141 1560
rect -175 1526 -141 1556
rect -17 2610 17 2640
rect -17 2606 17 2610
rect -17 2542 17 2568
rect -17 2534 17 2542
rect -17 2474 17 2496
rect -17 2462 17 2474
rect -17 2406 17 2424
rect -17 2390 17 2406
rect -17 2338 17 2352
rect -17 2318 17 2338
rect -17 2270 17 2280
rect -17 2246 17 2270
rect -17 2202 17 2208
rect -17 2174 17 2202
rect -17 2134 17 2136
rect -17 2102 17 2134
rect -17 2032 17 2064
rect -17 2030 17 2032
rect -17 1964 17 1992
rect -17 1958 17 1964
rect -17 1896 17 1920
rect -17 1886 17 1896
rect -17 1828 17 1848
rect -17 1814 17 1828
rect -17 1760 17 1776
rect -17 1742 17 1760
rect -17 1692 17 1704
rect -17 1670 17 1692
rect -17 1624 17 1632
rect -17 1598 17 1624
rect -17 1556 17 1560
rect -17 1526 17 1556
rect 141 2610 175 2640
rect 141 2606 175 2610
rect 141 2542 175 2568
rect 141 2534 175 2542
rect 141 2474 175 2496
rect 141 2462 175 2474
rect 141 2406 175 2424
rect 141 2390 175 2406
rect 141 2338 175 2352
rect 141 2318 175 2338
rect 141 2270 175 2280
rect 141 2246 175 2270
rect 141 2202 175 2208
rect 141 2174 175 2202
rect 141 2134 175 2136
rect 141 2102 175 2134
rect 141 2032 175 2064
rect 141 2030 175 2032
rect 141 1964 175 1992
rect 141 1958 175 1964
rect 141 1896 175 1920
rect 141 1886 175 1896
rect 141 1828 175 1848
rect 141 1814 175 1828
rect 141 1760 175 1776
rect 141 1742 175 1760
rect 141 1692 175 1704
rect 141 1670 175 1692
rect 141 1624 175 1632
rect 141 1598 175 1624
rect 141 1556 175 1560
rect 141 1526 175 1556
rect 299 2610 333 2640
rect 299 2606 333 2610
rect 299 2542 333 2568
rect 299 2534 333 2542
rect 299 2474 333 2496
rect 299 2462 333 2474
rect 299 2406 333 2424
rect 299 2390 333 2406
rect 299 2338 333 2352
rect 299 2318 333 2338
rect 299 2270 333 2280
rect 299 2246 333 2270
rect 299 2202 333 2208
rect 299 2174 333 2202
rect 299 2134 333 2136
rect 299 2102 333 2134
rect 299 2032 333 2064
rect 299 2030 333 2032
rect 299 1964 333 1992
rect 299 1958 333 1964
rect 299 1896 333 1920
rect 299 1886 333 1896
rect 299 1828 333 1848
rect 299 1814 333 1828
rect 299 1760 333 1776
rect 299 1742 333 1760
rect 299 1692 333 1704
rect 299 1670 333 1692
rect 299 1624 333 1632
rect 299 1598 333 1624
rect 299 1556 333 1560
rect 299 1526 333 1556
rect 457 2610 491 2640
rect 457 2606 491 2610
rect 457 2542 491 2568
rect 457 2534 491 2542
rect 457 2474 491 2496
rect 457 2462 491 2474
rect 457 2406 491 2424
rect 457 2390 491 2406
rect 457 2338 491 2352
rect 457 2318 491 2338
rect 457 2270 491 2280
rect 457 2246 491 2270
rect 457 2202 491 2208
rect 457 2174 491 2202
rect 457 2134 491 2136
rect 457 2102 491 2134
rect 457 2032 491 2064
rect 457 2030 491 2032
rect 457 1964 491 1992
rect 457 1958 491 1964
rect 457 1896 491 1920
rect 457 1886 491 1896
rect 457 1828 491 1848
rect 457 1814 491 1828
rect 457 1760 491 1776
rect 457 1742 491 1760
rect 457 1692 491 1704
rect 457 1670 491 1692
rect 457 1624 491 1632
rect 457 1598 491 1624
rect 457 1556 491 1560
rect 457 1526 491 1556
rect 615 2610 649 2640
rect 615 2606 649 2610
rect 615 2542 649 2568
rect 615 2534 649 2542
rect 615 2474 649 2496
rect 615 2462 649 2474
rect 615 2406 649 2424
rect 615 2390 649 2406
rect 615 2338 649 2352
rect 615 2318 649 2338
rect 615 2270 649 2280
rect 615 2246 649 2270
rect 615 2202 649 2208
rect 615 2174 649 2202
rect 615 2134 649 2136
rect 615 2102 649 2134
rect 615 2032 649 2064
rect 615 2030 649 2032
rect 615 1964 649 1992
rect 615 1958 649 1964
rect 615 1896 649 1920
rect 615 1886 649 1896
rect 615 1828 649 1848
rect 615 1814 649 1828
rect 615 1760 649 1776
rect 615 1742 649 1760
rect 615 1692 649 1704
rect 615 1670 649 1692
rect 615 1624 649 1632
rect 615 1598 649 1624
rect 615 1556 649 1560
rect 615 1526 649 1556
rect 773 2610 807 2640
rect 773 2606 807 2610
rect 773 2542 807 2568
rect 773 2534 807 2542
rect 773 2474 807 2496
rect 773 2462 807 2474
rect 773 2406 807 2424
rect 773 2390 807 2406
rect 773 2338 807 2352
rect 773 2318 807 2338
rect 773 2270 807 2280
rect 773 2246 807 2270
rect 773 2202 807 2208
rect 773 2174 807 2202
rect 773 2134 807 2136
rect 773 2102 807 2134
rect 773 2032 807 2064
rect 773 2030 807 2032
rect 773 1964 807 1992
rect 773 1958 807 1964
rect 773 1896 807 1920
rect 773 1886 807 1896
rect 773 1828 807 1848
rect 773 1814 807 1828
rect 773 1760 807 1776
rect 773 1742 807 1760
rect 773 1692 807 1704
rect 773 1670 807 1692
rect 773 1624 807 1632
rect 773 1598 807 1624
rect 773 1556 807 1560
rect 773 1526 807 1556
rect 931 2610 965 2640
rect 931 2606 965 2610
rect 931 2542 965 2568
rect 931 2534 965 2542
rect 931 2474 965 2496
rect 931 2462 965 2474
rect 931 2406 965 2424
rect 931 2390 965 2406
rect 931 2338 965 2352
rect 931 2318 965 2338
rect 931 2270 965 2280
rect 931 2246 965 2270
rect 931 2202 965 2208
rect 931 2174 965 2202
rect 931 2134 965 2136
rect 931 2102 965 2134
rect 931 2032 965 2064
rect 931 2030 965 2032
rect 931 1964 965 1992
rect 931 1958 965 1964
rect 931 1896 965 1920
rect 931 1886 965 1896
rect 931 1828 965 1848
rect 931 1814 965 1828
rect 931 1760 965 1776
rect 931 1742 965 1760
rect 931 1692 965 1704
rect 931 1670 965 1692
rect 931 1624 965 1632
rect 931 1598 965 1624
rect 931 1556 965 1560
rect 931 1526 965 1556
rect 1089 2610 1123 2640
rect 1089 2606 1123 2610
rect 1089 2542 1123 2568
rect 1089 2534 1123 2542
rect 1089 2474 1123 2496
rect 1089 2462 1123 2474
rect 1089 2406 1123 2424
rect 1089 2390 1123 2406
rect 1089 2338 1123 2352
rect 1089 2318 1123 2338
rect 1089 2270 1123 2280
rect 1089 2246 1123 2270
rect 1089 2202 1123 2208
rect 1089 2174 1123 2202
rect 1089 2134 1123 2136
rect 1089 2102 1123 2134
rect 1089 2032 1123 2064
rect 1089 2030 1123 2032
rect 1089 1964 1123 1992
rect 1089 1958 1123 1964
rect 1089 1896 1123 1920
rect 1089 1886 1123 1896
rect 1089 1828 1123 1848
rect 1089 1814 1123 1828
rect 1089 1760 1123 1776
rect 1089 1742 1123 1760
rect 1089 1692 1123 1704
rect 1089 1670 1123 1692
rect 1089 1624 1123 1632
rect 1089 1598 1123 1624
rect 1089 1556 1123 1560
rect 1089 1526 1123 1556
rect -1044 1402 -1010 1436
rect -886 1402 -852 1436
rect -728 1402 -694 1436
rect -570 1402 -536 1436
rect -412 1402 -378 1436
rect -254 1402 -220 1436
rect -96 1402 -62 1436
rect 62 1402 96 1436
rect 220 1402 254 1436
rect 378 1402 412 1436
rect 536 1402 570 1436
rect 694 1402 728 1436
rect 852 1402 886 1436
rect 1010 1402 1044 1436
rect -1123 1245 -1089 1275
rect -1123 1241 -1089 1245
rect -1123 1177 -1089 1203
rect -1123 1169 -1089 1177
rect -1123 1109 -1089 1131
rect -1123 1097 -1089 1109
rect -1123 1041 -1089 1059
rect -1123 1025 -1089 1041
rect -1123 973 -1089 987
rect -1123 953 -1089 973
rect -1123 905 -1089 915
rect -1123 881 -1089 905
rect -1123 837 -1089 843
rect -1123 809 -1089 837
rect -1123 769 -1089 771
rect -1123 737 -1089 769
rect -1123 667 -1089 699
rect -1123 665 -1089 667
rect -1123 599 -1089 627
rect -1123 593 -1089 599
rect -1123 531 -1089 555
rect -1123 521 -1089 531
rect -1123 463 -1089 483
rect -1123 449 -1089 463
rect -1123 395 -1089 411
rect -1123 377 -1089 395
rect -1123 327 -1089 339
rect -1123 305 -1089 327
rect -1123 259 -1089 267
rect -1123 233 -1089 259
rect -1123 191 -1089 195
rect -1123 161 -1089 191
rect -965 1245 -931 1275
rect -965 1241 -931 1245
rect -965 1177 -931 1203
rect -965 1169 -931 1177
rect -965 1109 -931 1131
rect -965 1097 -931 1109
rect -965 1041 -931 1059
rect -965 1025 -931 1041
rect -965 973 -931 987
rect -965 953 -931 973
rect -965 905 -931 915
rect -965 881 -931 905
rect -965 837 -931 843
rect -965 809 -931 837
rect -965 769 -931 771
rect -965 737 -931 769
rect -965 667 -931 699
rect -965 665 -931 667
rect -965 599 -931 627
rect -965 593 -931 599
rect -965 531 -931 555
rect -965 521 -931 531
rect -965 463 -931 483
rect -965 449 -931 463
rect -965 395 -931 411
rect -965 377 -931 395
rect -965 327 -931 339
rect -965 305 -931 327
rect -965 259 -931 267
rect -965 233 -931 259
rect -965 191 -931 195
rect -965 161 -931 191
rect -807 1245 -773 1275
rect -807 1241 -773 1245
rect -807 1177 -773 1203
rect -807 1169 -773 1177
rect -807 1109 -773 1131
rect -807 1097 -773 1109
rect -807 1041 -773 1059
rect -807 1025 -773 1041
rect -807 973 -773 987
rect -807 953 -773 973
rect -807 905 -773 915
rect -807 881 -773 905
rect -807 837 -773 843
rect -807 809 -773 837
rect -807 769 -773 771
rect -807 737 -773 769
rect -807 667 -773 699
rect -807 665 -773 667
rect -807 599 -773 627
rect -807 593 -773 599
rect -807 531 -773 555
rect -807 521 -773 531
rect -807 463 -773 483
rect -807 449 -773 463
rect -807 395 -773 411
rect -807 377 -773 395
rect -807 327 -773 339
rect -807 305 -773 327
rect -807 259 -773 267
rect -807 233 -773 259
rect -807 191 -773 195
rect -807 161 -773 191
rect -649 1245 -615 1275
rect -649 1241 -615 1245
rect -649 1177 -615 1203
rect -649 1169 -615 1177
rect -649 1109 -615 1131
rect -649 1097 -615 1109
rect -649 1041 -615 1059
rect -649 1025 -615 1041
rect -649 973 -615 987
rect -649 953 -615 973
rect -649 905 -615 915
rect -649 881 -615 905
rect -649 837 -615 843
rect -649 809 -615 837
rect -649 769 -615 771
rect -649 737 -615 769
rect -649 667 -615 699
rect -649 665 -615 667
rect -649 599 -615 627
rect -649 593 -615 599
rect -649 531 -615 555
rect -649 521 -615 531
rect -649 463 -615 483
rect -649 449 -615 463
rect -649 395 -615 411
rect -649 377 -615 395
rect -649 327 -615 339
rect -649 305 -615 327
rect -649 259 -615 267
rect -649 233 -615 259
rect -649 191 -615 195
rect -649 161 -615 191
rect -491 1245 -457 1275
rect -491 1241 -457 1245
rect -491 1177 -457 1203
rect -491 1169 -457 1177
rect -491 1109 -457 1131
rect -491 1097 -457 1109
rect -491 1041 -457 1059
rect -491 1025 -457 1041
rect -491 973 -457 987
rect -491 953 -457 973
rect -491 905 -457 915
rect -491 881 -457 905
rect -491 837 -457 843
rect -491 809 -457 837
rect -491 769 -457 771
rect -491 737 -457 769
rect -491 667 -457 699
rect -491 665 -457 667
rect -491 599 -457 627
rect -491 593 -457 599
rect -491 531 -457 555
rect -491 521 -457 531
rect -491 463 -457 483
rect -491 449 -457 463
rect -491 395 -457 411
rect -491 377 -457 395
rect -491 327 -457 339
rect -491 305 -457 327
rect -491 259 -457 267
rect -491 233 -457 259
rect -491 191 -457 195
rect -491 161 -457 191
rect -333 1245 -299 1275
rect -333 1241 -299 1245
rect -333 1177 -299 1203
rect -333 1169 -299 1177
rect -333 1109 -299 1131
rect -333 1097 -299 1109
rect -333 1041 -299 1059
rect -333 1025 -299 1041
rect -333 973 -299 987
rect -333 953 -299 973
rect -333 905 -299 915
rect -333 881 -299 905
rect -333 837 -299 843
rect -333 809 -299 837
rect -333 769 -299 771
rect -333 737 -299 769
rect -333 667 -299 699
rect -333 665 -299 667
rect -333 599 -299 627
rect -333 593 -299 599
rect -333 531 -299 555
rect -333 521 -299 531
rect -333 463 -299 483
rect -333 449 -299 463
rect -333 395 -299 411
rect -333 377 -299 395
rect -333 327 -299 339
rect -333 305 -299 327
rect -333 259 -299 267
rect -333 233 -299 259
rect -333 191 -299 195
rect -333 161 -299 191
rect -175 1245 -141 1275
rect -175 1241 -141 1245
rect -175 1177 -141 1203
rect -175 1169 -141 1177
rect -175 1109 -141 1131
rect -175 1097 -141 1109
rect -175 1041 -141 1059
rect -175 1025 -141 1041
rect -175 973 -141 987
rect -175 953 -141 973
rect -175 905 -141 915
rect -175 881 -141 905
rect -175 837 -141 843
rect -175 809 -141 837
rect -175 769 -141 771
rect -175 737 -141 769
rect -175 667 -141 699
rect -175 665 -141 667
rect -175 599 -141 627
rect -175 593 -141 599
rect -175 531 -141 555
rect -175 521 -141 531
rect -175 463 -141 483
rect -175 449 -141 463
rect -175 395 -141 411
rect -175 377 -141 395
rect -175 327 -141 339
rect -175 305 -141 327
rect -175 259 -141 267
rect -175 233 -141 259
rect -175 191 -141 195
rect -175 161 -141 191
rect -17 1245 17 1275
rect -17 1241 17 1245
rect -17 1177 17 1203
rect -17 1169 17 1177
rect -17 1109 17 1131
rect -17 1097 17 1109
rect -17 1041 17 1059
rect -17 1025 17 1041
rect -17 973 17 987
rect -17 953 17 973
rect -17 905 17 915
rect -17 881 17 905
rect -17 837 17 843
rect -17 809 17 837
rect -17 769 17 771
rect -17 737 17 769
rect -17 667 17 699
rect -17 665 17 667
rect -17 599 17 627
rect -17 593 17 599
rect -17 531 17 555
rect -17 521 17 531
rect -17 463 17 483
rect -17 449 17 463
rect -17 395 17 411
rect -17 377 17 395
rect -17 327 17 339
rect -17 305 17 327
rect -17 259 17 267
rect -17 233 17 259
rect -17 191 17 195
rect -17 161 17 191
rect 141 1245 175 1275
rect 141 1241 175 1245
rect 141 1177 175 1203
rect 141 1169 175 1177
rect 141 1109 175 1131
rect 141 1097 175 1109
rect 141 1041 175 1059
rect 141 1025 175 1041
rect 141 973 175 987
rect 141 953 175 973
rect 141 905 175 915
rect 141 881 175 905
rect 141 837 175 843
rect 141 809 175 837
rect 141 769 175 771
rect 141 737 175 769
rect 141 667 175 699
rect 141 665 175 667
rect 141 599 175 627
rect 141 593 175 599
rect 141 531 175 555
rect 141 521 175 531
rect 141 463 175 483
rect 141 449 175 463
rect 141 395 175 411
rect 141 377 175 395
rect 141 327 175 339
rect 141 305 175 327
rect 141 259 175 267
rect 141 233 175 259
rect 141 191 175 195
rect 141 161 175 191
rect 299 1245 333 1275
rect 299 1241 333 1245
rect 299 1177 333 1203
rect 299 1169 333 1177
rect 299 1109 333 1131
rect 299 1097 333 1109
rect 299 1041 333 1059
rect 299 1025 333 1041
rect 299 973 333 987
rect 299 953 333 973
rect 299 905 333 915
rect 299 881 333 905
rect 299 837 333 843
rect 299 809 333 837
rect 299 769 333 771
rect 299 737 333 769
rect 299 667 333 699
rect 299 665 333 667
rect 299 599 333 627
rect 299 593 333 599
rect 299 531 333 555
rect 299 521 333 531
rect 299 463 333 483
rect 299 449 333 463
rect 299 395 333 411
rect 299 377 333 395
rect 299 327 333 339
rect 299 305 333 327
rect 299 259 333 267
rect 299 233 333 259
rect 299 191 333 195
rect 299 161 333 191
rect 457 1245 491 1275
rect 457 1241 491 1245
rect 457 1177 491 1203
rect 457 1169 491 1177
rect 457 1109 491 1131
rect 457 1097 491 1109
rect 457 1041 491 1059
rect 457 1025 491 1041
rect 457 973 491 987
rect 457 953 491 973
rect 457 905 491 915
rect 457 881 491 905
rect 457 837 491 843
rect 457 809 491 837
rect 457 769 491 771
rect 457 737 491 769
rect 457 667 491 699
rect 457 665 491 667
rect 457 599 491 627
rect 457 593 491 599
rect 457 531 491 555
rect 457 521 491 531
rect 457 463 491 483
rect 457 449 491 463
rect 457 395 491 411
rect 457 377 491 395
rect 457 327 491 339
rect 457 305 491 327
rect 457 259 491 267
rect 457 233 491 259
rect 457 191 491 195
rect 457 161 491 191
rect 615 1245 649 1275
rect 615 1241 649 1245
rect 615 1177 649 1203
rect 615 1169 649 1177
rect 615 1109 649 1131
rect 615 1097 649 1109
rect 615 1041 649 1059
rect 615 1025 649 1041
rect 615 973 649 987
rect 615 953 649 973
rect 615 905 649 915
rect 615 881 649 905
rect 615 837 649 843
rect 615 809 649 837
rect 615 769 649 771
rect 615 737 649 769
rect 615 667 649 699
rect 615 665 649 667
rect 615 599 649 627
rect 615 593 649 599
rect 615 531 649 555
rect 615 521 649 531
rect 615 463 649 483
rect 615 449 649 463
rect 615 395 649 411
rect 615 377 649 395
rect 615 327 649 339
rect 615 305 649 327
rect 615 259 649 267
rect 615 233 649 259
rect 615 191 649 195
rect 615 161 649 191
rect 773 1245 807 1275
rect 773 1241 807 1245
rect 773 1177 807 1203
rect 773 1169 807 1177
rect 773 1109 807 1131
rect 773 1097 807 1109
rect 773 1041 807 1059
rect 773 1025 807 1041
rect 773 973 807 987
rect 773 953 807 973
rect 773 905 807 915
rect 773 881 807 905
rect 773 837 807 843
rect 773 809 807 837
rect 773 769 807 771
rect 773 737 807 769
rect 773 667 807 699
rect 773 665 807 667
rect 773 599 807 627
rect 773 593 807 599
rect 773 531 807 555
rect 773 521 807 531
rect 773 463 807 483
rect 773 449 807 463
rect 773 395 807 411
rect 773 377 807 395
rect 773 327 807 339
rect 773 305 807 327
rect 773 259 807 267
rect 773 233 807 259
rect 773 191 807 195
rect 773 161 807 191
rect 931 1245 965 1275
rect 931 1241 965 1245
rect 931 1177 965 1203
rect 931 1169 965 1177
rect 931 1109 965 1131
rect 931 1097 965 1109
rect 931 1041 965 1059
rect 931 1025 965 1041
rect 931 973 965 987
rect 931 953 965 973
rect 931 905 965 915
rect 931 881 965 905
rect 931 837 965 843
rect 931 809 965 837
rect 931 769 965 771
rect 931 737 965 769
rect 931 667 965 699
rect 931 665 965 667
rect 931 599 965 627
rect 931 593 965 599
rect 931 531 965 555
rect 931 521 965 531
rect 931 463 965 483
rect 931 449 965 463
rect 931 395 965 411
rect 931 377 965 395
rect 931 327 965 339
rect 931 305 965 327
rect 931 259 965 267
rect 931 233 965 259
rect 931 191 965 195
rect 931 161 965 191
rect 1089 1245 1123 1275
rect 1089 1241 1123 1245
rect 1089 1177 1123 1203
rect 1089 1169 1123 1177
rect 1089 1109 1123 1131
rect 1089 1097 1123 1109
rect 1089 1041 1123 1059
rect 1089 1025 1123 1041
rect 1089 973 1123 987
rect 1089 953 1123 973
rect 1089 905 1123 915
rect 1089 881 1123 905
rect 1089 837 1123 843
rect 1089 809 1123 837
rect 1089 769 1123 771
rect 1089 737 1123 769
rect 1089 667 1123 699
rect 1089 665 1123 667
rect 1089 599 1123 627
rect 1089 593 1123 599
rect 1089 531 1123 555
rect 1089 521 1123 531
rect 1089 463 1123 483
rect 1089 449 1123 463
rect 1089 395 1123 411
rect 1089 377 1123 395
rect 1089 327 1123 339
rect 1089 305 1123 327
rect 1089 259 1123 267
rect 1089 233 1123 259
rect 1089 191 1123 195
rect 1089 161 1123 191
rect -1044 37 -1010 71
rect -886 37 -852 71
rect -728 37 -694 71
rect -570 37 -536 71
rect -412 37 -378 71
rect -254 37 -220 71
rect -96 37 -62 71
rect 62 37 96 71
rect 220 37 254 71
rect 378 37 412 71
rect 536 37 570 71
rect 694 37 728 71
rect 852 37 886 71
rect 1010 37 1044 71
rect -1123 -120 -1089 -90
rect -1123 -124 -1089 -120
rect -1123 -188 -1089 -162
rect -1123 -196 -1089 -188
rect -1123 -256 -1089 -234
rect -1123 -268 -1089 -256
rect -1123 -324 -1089 -306
rect -1123 -340 -1089 -324
rect -1123 -392 -1089 -378
rect -1123 -412 -1089 -392
rect -1123 -460 -1089 -450
rect -1123 -484 -1089 -460
rect -1123 -528 -1089 -522
rect -1123 -556 -1089 -528
rect -1123 -596 -1089 -594
rect -1123 -628 -1089 -596
rect -1123 -698 -1089 -666
rect -1123 -700 -1089 -698
rect -1123 -766 -1089 -738
rect -1123 -772 -1089 -766
rect -1123 -834 -1089 -810
rect -1123 -844 -1089 -834
rect -1123 -902 -1089 -882
rect -1123 -916 -1089 -902
rect -1123 -970 -1089 -954
rect -1123 -988 -1089 -970
rect -1123 -1038 -1089 -1026
rect -1123 -1060 -1089 -1038
rect -1123 -1106 -1089 -1098
rect -1123 -1132 -1089 -1106
rect -1123 -1174 -1089 -1170
rect -1123 -1204 -1089 -1174
rect -965 -120 -931 -90
rect -965 -124 -931 -120
rect -965 -188 -931 -162
rect -965 -196 -931 -188
rect -965 -256 -931 -234
rect -965 -268 -931 -256
rect -965 -324 -931 -306
rect -965 -340 -931 -324
rect -965 -392 -931 -378
rect -965 -412 -931 -392
rect -965 -460 -931 -450
rect -965 -484 -931 -460
rect -965 -528 -931 -522
rect -965 -556 -931 -528
rect -965 -596 -931 -594
rect -965 -628 -931 -596
rect -965 -698 -931 -666
rect -965 -700 -931 -698
rect -965 -766 -931 -738
rect -965 -772 -931 -766
rect -965 -834 -931 -810
rect -965 -844 -931 -834
rect -965 -902 -931 -882
rect -965 -916 -931 -902
rect -965 -970 -931 -954
rect -965 -988 -931 -970
rect -965 -1038 -931 -1026
rect -965 -1060 -931 -1038
rect -965 -1106 -931 -1098
rect -965 -1132 -931 -1106
rect -965 -1174 -931 -1170
rect -965 -1204 -931 -1174
rect -807 -120 -773 -90
rect -807 -124 -773 -120
rect -807 -188 -773 -162
rect -807 -196 -773 -188
rect -807 -256 -773 -234
rect -807 -268 -773 -256
rect -807 -324 -773 -306
rect -807 -340 -773 -324
rect -807 -392 -773 -378
rect -807 -412 -773 -392
rect -807 -460 -773 -450
rect -807 -484 -773 -460
rect -807 -528 -773 -522
rect -807 -556 -773 -528
rect -807 -596 -773 -594
rect -807 -628 -773 -596
rect -807 -698 -773 -666
rect -807 -700 -773 -698
rect -807 -766 -773 -738
rect -807 -772 -773 -766
rect -807 -834 -773 -810
rect -807 -844 -773 -834
rect -807 -902 -773 -882
rect -807 -916 -773 -902
rect -807 -970 -773 -954
rect -807 -988 -773 -970
rect -807 -1038 -773 -1026
rect -807 -1060 -773 -1038
rect -807 -1106 -773 -1098
rect -807 -1132 -773 -1106
rect -807 -1174 -773 -1170
rect -807 -1204 -773 -1174
rect -649 -120 -615 -90
rect -649 -124 -615 -120
rect -649 -188 -615 -162
rect -649 -196 -615 -188
rect -649 -256 -615 -234
rect -649 -268 -615 -256
rect -649 -324 -615 -306
rect -649 -340 -615 -324
rect -649 -392 -615 -378
rect -649 -412 -615 -392
rect -649 -460 -615 -450
rect -649 -484 -615 -460
rect -649 -528 -615 -522
rect -649 -556 -615 -528
rect -649 -596 -615 -594
rect -649 -628 -615 -596
rect -649 -698 -615 -666
rect -649 -700 -615 -698
rect -649 -766 -615 -738
rect -649 -772 -615 -766
rect -649 -834 -615 -810
rect -649 -844 -615 -834
rect -649 -902 -615 -882
rect -649 -916 -615 -902
rect -649 -970 -615 -954
rect -649 -988 -615 -970
rect -649 -1038 -615 -1026
rect -649 -1060 -615 -1038
rect -649 -1106 -615 -1098
rect -649 -1132 -615 -1106
rect -649 -1174 -615 -1170
rect -649 -1204 -615 -1174
rect -491 -120 -457 -90
rect -491 -124 -457 -120
rect -491 -188 -457 -162
rect -491 -196 -457 -188
rect -491 -256 -457 -234
rect -491 -268 -457 -256
rect -491 -324 -457 -306
rect -491 -340 -457 -324
rect -491 -392 -457 -378
rect -491 -412 -457 -392
rect -491 -460 -457 -450
rect -491 -484 -457 -460
rect -491 -528 -457 -522
rect -491 -556 -457 -528
rect -491 -596 -457 -594
rect -491 -628 -457 -596
rect -491 -698 -457 -666
rect -491 -700 -457 -698
rect -491 -766 -457 -738
rect -491 -772 -457 -766
rect -491 -834 -457 -810
rect -491 -844 -457 -834
rect -491 -902 -457 -882
rect -491 -916 -457 -902
rect -491 -970 -457 -954
rect -491 -988 -457 -970
rect -491 -1038 -457 -1026
rect -491 -1060 -457 -1038
rect -491 -1106 -457 -1098
rect -491 -1132 -457 -1106
rect -491 -1174 -457 -1170
rect -491 -1204 -457 -1174
rect -333 -120 -299 -90
rect -333 -124 -299 -120
rect -333 -188 -299 -162
rect -333 -196 -299 -188
rect -333 -256 -299 -234
rect -333 -268 -299 -256
rect -333 -324 -299 -306
rect -333 -340 -299 -324
rect -333 -392 -299 -378
rect -333 -412 -299 -392
rect -333 -460 -299 -450
rect -333 -484 -299 -460
rect -333 -528 -299 -522
rect -333 -556 -299 -528
rect -333 -596 -299 -594
rect -333 -628 -299 -596
rect -333 -698 -299 -666
rect -333 -700 -299 -698
rect -333 -766 -299 -738
rect -333 -772 -299 -766
rect -333 -834 -299 -810
rect -333 -844 -299 -834
rect -333 -902 -299 -882
rect -333 -916 -299 -902
rect -333 -970 -299 -954
rect -333 -988 -299 -970
rect -333 -1038 -299 -1026
rect -333 -1060 -299 -1038
rect -333 -1106 -299 -1098
rect -333 -1132 -299 -1106
rect -333 -1174 -299 -1170
rect -333 -1204 -299 -1174
rect -175 -120 -141 -90
rect -175 -124 -141 -120
rect -175 -188 -141 -162
rect -175 -196 -141 -188
rect -175 -256 -141 -234
rect -175 -268 -141 -256
rect -175 -324 -141 -306
rect -175 -340 -141 -324
rect -175 -392 -141 -378
rect -175 -412 -141 -392
rect -175 -460 -141 -450
rect -175 -484 -141 -460
rect -175 -528 -141 -522
rect -175 -556 -141 -528
rect -175 -596 -141 -594
rect -175 -628 -141 -596
rect -175 -698 -141 -666
rect -175 -700 -141 -698
rect -175 -766 -141 -738
rect -175 -772 -141 -766
rect -175 -834 -141 -810
rect -175 -844 -141 -834
rect -175 -902 -141 -882
rect -175 -916 -141 -902
rect -175 -970 -141 -954
rect -175 -988 -141 -970
rect -175 -1038 -141 -1026
rect -175 -1060 -141 -1038
rect -175 -1106 -141 -1098
rect -175 -1132 -141 -1106
rect -175 -1174 -141 -1170
rect -175 -1204 -141 -1174
rect -17 -120 17 -90
rect -17 -124 17 -120
rect -17 -188 17 -162
rect -17 -196 17 -188
rect -17 -256 17 -234
rect -17 -268 17 -256
rect -17 -324 17 -306
rect -17 -340 17 -324
rect -17 -392 17 -378
rect -17 -412 17 -392
rect -17 -460 17 -450
rect -17 -484 17 -460
rect -17 -528 17 -522
rect -17 -556 17 -528
rect -17 -596 17 -594
rect -17 -628 17 -596
rect -17 -698 17 -666
rect -17 -700 17 -698
rect -17 -766 17 -738
rect -17 -772 17 -766
rect -17 -834 17 -810
rect -17 -844 17 -834
rect -17 -902 17 -882
rect -17 -916 17 -902
rect -17 -970 17 -954
rect -17 -988 17 -970
rect -17 -1038 17 -1026
rect -17 -1060 17 -1038
rect -17 -1106 17 -1098
rect -17 -1132 17 -1106
rect -17 -1174 17 -1170
rect -17 -1204 17 -1174
rect 141 -120 175 -90
rect 141 -124 175 -120
rect 141 -188 175 -162
rect 141 -196 175 -188
rect 141 -256 175 -234
rect 141 -268 175 -256
rect 141 -324 175 -306
rect 141 -340 175 -324
rect 141 -392 175 -378
rect 141 -412 175 -392
rect 141 -460 175 -450
rect 141 -484 175 -460
rect 141 -528 175 -522
rect 141 -556 175 -528
rect 141 -596 175 -594
rect 141 -628 175 -596
rect 141 -698 175 -666
rect 141 -700 175 -698
rect 141 -766 175 -738
rect 141 -772 175 -766
rect 141 -834 175 -810
rect 141 -844 175 -834
rect 141 -902 175 -882
rect 141 -916 175 -902
rect 141 -970 175 -954
rect 141 -988 175 -970
rect 141 -1038 175 -1026
rect 141 -1060 175 -1038
rect 141 -1106 175 -1098
rect 141 -1132 175 -1106
rect 141 -1174 175 -1170
rect 141 -1204 175 -1174
rect 299 -120 333 -90
rect 299 -124 333 -120
rect 299 -188 333 -162
rect 299 -196 333 -188
rect 299 -256 333 -234
rect 299 -268 333 -256
rect 299 -324 333 -306
rect 299 -340 333 -324
rect 299 -392 333 -378
rect 299 -412 333 -392
rect 299 -460 333 -450
rect 299 -484 333 -460
rect 299 -528 333 -522
rect 299 -556 333 -528
rect 299 -596 333 -594
rect 299 -628 333 -596
rect 299 -698 333 -666
rect 299 -700 333 -698
rect 299 -766 333 -738
rect 299 -772 333 -766
rect 299 -834 333 -810
rect 299 -844 333 -834
rect 299 -902 333 -882
rect 299 -916 333 -902
rect 299 -970 333 -954
rect 299 -988 333 -970
rect 299 -1038 333 -1026
rect 299 -1060 333 -1038
rect 299 -1106 333 -1098
rect 299 -1132 333 -1106
rect 299 -1174 333 -1170
rect 299 -1204 333 -1174
rect 457 -120 491 -90
rect 457 -124 491 -120
rect 457 -188 491 -162
rect 457 -196 491 -188
rect 457 -256 491 -234
rect 457 -268 491 -256
rect 457 -324 491 -306
rect 457 -340 491 -324
rect 457 -392 491 -378
rect 457 -412 491 -392
rect 457 -460 491 -450
rect 457 -484 491 -460
rect 457 -528 491 -522
rect 457 -556 491 -528
rect 457 -596 491 -594
rect 457 -628 491 -596
rect 457 -698 491 -666
rect 457 -700 491 -698
rect 457 -766 491 -738
rect 457 -772 491 -766
rect 457 -834 491 -810
rect 457 -844 491 -834
rect 457 -902 491 -882
rect 457 -916 491 -902
rect 457 -970 491 -954
rect 457 -988 491 -970
rect 457 -1038 491 -1026
rect 457 -1060 491 -1038
rect 457 -1106 491 -1098
rect 457 -1132 491 -1106
rect 457 -1174 491 -1170
rect 457 -1204 491 -1174
rect 615 -120 649 -90
rect 615 -124 649 -120
rect 615 -188 649 -162
rect 615 -196 649 -188
rect 615 -256 649 -234
rect 615 -268 649 -256
rect 615 -324 649 -306
rect 615 -340 649 -324
rect 615 -392 649 -378
rect 615 -412 649 -392
rect 615 -460 649 -450
rect 615 -484 649 -460
rect 615 -528 649 -522
rect 615 -556 649 -528
rect 615 -596 649 -594
rect 615 -628 649 -596
rect 615 -698 649 -666
rect 615 -700 649 -698
rect 615 -766 649 -738
rect 615 -772 649 -766
rect 615 -834 649 -810
rect 615 -844 649 -834
rect 615 -902 649 -882
rect 615 -916 649 -902
rect 615 -970 649 -954
rect 615 -988 649 -970
rect 615 -1038 649 -1026
rect 615 -1060 649 -1038
rect 615 -1106 649 -1098
rect 615 -1132 649 -1106
rect 615 -1174 649 -1170
rect 615 -1204 649 -1174
rect 773 -120 807 -90
rect 773 -124 807 -120
rect 773 -188 807 -162
rect 773 -196 807 -188
rect 773 -256 807 -234
rect 773 -268 807 -256
rect 773 -324 807 -306
rect 773 -340 807 -324
rect 773 -392 807 -378
rect 773 -412 807 -392
rect 773 -460 807 -450
rect 773 -484 807 -460
rect 773 -528 807 -522
rect 773 -556 807 -528
rect 773 -596 807 -594
rect 773 -628 807 -596
rect 773 -698 807 -666
rect 773 -700 807 -698
rect 773 -766 807 -738
rect 773 -772 807 -766
rect 773 -834 807 -810
rect 773 -844 807 -834
rect 773 -902 807 -882
rect 773 -916 807 -902
rect 773 -970 807 -954
rect 773 -988 807 -970
rect 773 -1038 807 -1026
rect 773 -1060 807 -1038
rect 773 -1106 807 -1098
rect 773 -1132 807 -1106
rect 773 -1174 807 -1170
rect 773 -1204 807 -1174
rect 931 -120 965 -90
rect 931 -124 965 -120
rect 931 -188 965 -162
rect 931 -196 965 -188
rect 931 -256 965 -234
rect 931 -268 965 -256
rect 931 -324 965 -306
rect 931 -340 965 -324
rect 931 -392 965 -378
rect 931 -412 965 -392
rect 931 -460 965 -450
rect 931 -484 965 -460
rect 931 -528 965 -522
rect 931 -556 965 -528
rect 931 -596 965 -594
rect 931 -628 965 -596
rect 931 -698 965 -666
rect 931 -700 965 -698
rect 931 -766 965 -738
rect 931 -772 965 -766
rect 931 -834 965 -810
rect 931 -844 965 -834
rect 931 -902 965 -882
rect 931 -916 965 -902
rect 931 -970 965 -954
rect 931 -988 965 -970
rect 931 -1038 965 -1026
rect 931 -1060 965 -1038
rect 931 -1106 965 -1098
rect 931 -1132 965 -1106
rect 931 -1174 965 -1170
rect 931 -1204 965 -1174
rect 1089 -120 1123 -90
rect 1089 -124 1123 -120
rect 1089 -188 1123 -162
rect 1089 -196 1123 -188
rect 1089 -256 1123 -234
rect 1089 -268 1123 -256
rect 1089 -324 1123 -306
rect 1089 -340 1123 -324
rect 1089 -392 1123 -378
rect 1089 -412 1123 -392
rect 1089 -460 1123 -450
rect 1089 -484 1123 -460
rect 1089 -528 1123 -522
rect 1089 -556 1123 -528
rect 1089 -596 1123 -594
rect 1089 -628 1123 -596
rect 1089 -698 1123 -666
rect 1089 -700 1123 -698
rect 1089 -766 1123 -738
rect 1089 -772 1123 -766
rect 1089 -834 1123 -810
rect 1089 -844 1123 -834
rect 1089 -902 1123 -882
rect 1089 -916 1123 -902
rect 1089 -970 1123 -954
rect 1089 -988 1123 -970
rect 1089 -1038 1123 -1026
rect 1089 -1060 1123 -1038
rect 1089 -1106 1123 -1098
rect 1089 -1132 1123 -1106
rect 1089 -1174 1123 -1170
rect 1089 -1204 1123 -1174
rect -1044 -1328 -1010 -1294
rect -886 -1328 -852 -1294
rect -728 -1328 -694 -1294
rect -570 -1328 -536 -1294
rect -412 -1328 -378 -1294
rect -254 -1328 -220 -1294
rect -96 -1328 -62 -1294
rect 62 -1328 96 -1294
rect 220 -1328 254 -1294
rect 378 -1328 412 -1294
rect 536 -1328 570 -1294
rect 694 -1328 728 -1294
rect 852 -1328 886 -1294
rect 1010 -1328 1044 -1294
rect -1123 -1485 -1089 -1455
rect -1123 -1489 -1089 -1485
rect -1123 -1553 -1089 -1527
rect -1123 -1561 -1089 -1553
rect -1123 -1621 -1089 -1599
rect -1123 -1633 -1089 -1621
rect -1123 -1689 -1089 -1671
rect -1123 -1705 -1089 -1689
rect -1123 -1757 -1089 -1743
rect -1123 -1777 -1089 -1757
rect -1123 -1825 -1089 -1815
rect -1123 -1849 -1089 -1825
rect -1123 -1893 -1089 -1887
rect -1123 -1921 -1089 -1893
rect -1123 -1961 -1089 -1959
rect -1123 -1993 -1089 -1961
rect -1123 -2063 -1089 -2031
rect -1123 -2065 -1089 -2063
rect -1123 -2131 -1089 -2103
rect -1123 -2137 -1089 -2131
rect -1123 -2199 -1089 -2175
rect -1123 -2209 -1089 -2199
rect -1123 -2267 -1089 -2247
rect -1123 -2281 -1089 -2267
rect -1123 -2335 -1089 -2319
rect -1123 -2353 -1089 -2335
rect -1123 -2403 -1089 -2391
rect -1123 -2425 -1089 -2403
rect -1123 -2471 -1089 -2463
rect -1123 -2497 -1089 -2471
rect -1123 -2539 -1089 -2535
rect -1123 -2569 -1089 -2539
rect -965 -1485 -931 -1455
rect -965 -1489 -931 -1485
rect -965 -1553 -931 -1527
rect -965 -1561 -931 -1553
rect -965 -1621 -931 -1599
rect -965 -1633 -931 -1621
rect -965 -1689 -931 -1671
rect -965 -1705 -931 -1689
rect -965 -1757 -931 -1743
rect -965 -1777 -931 -1757
rect -965 -1825 -931 -1815
rect -965 -1849 -931 -1825
rect -965 -1893 -931 -1887
rect -965 -1921 -931 -1893
rect -965 -1961 -931 -1959
rect -965 -1993 -931 -1961
rect -965 -2063 -931 -2031
rect -965 -2065 -931 -2063
rect -965 -2131 -931 -2103
rect -965 -2137 -931 -2131
rect -965 -2199 -931 -2175
rect -965 -2209 -931 -2199
rect -965 -2267 -931 -2247
rect -965 -2281 -931 -2267
rect -965 -2335 -931 -2319
rect -965 -2353 -931 -2335
rect -965 -2403 -931 -2391
rect -965 -2425 -931 -2403
rect -965 -2471 -931 -2463
rect -965 -2497 -931 -2471
rect -965 -2539 -931 -2535
rect -965 -2569 -931 -2539
rect -807 -1485 -773 -1455
rect -807 -1489 -773 -1485
rect -807 -1553 -773 -1527
rect -807 -1561 -773 -1553
rect -807 -1621 -773 -1599
rect -807 -1633 -773 -1621
rect -807 -1689 -773 -1671
rect -807 -1705 -773 -1689
rect -807 -1757 -773 -1743
rect -807 -1777 -773 -1757
rect -807 -1825 -773 -1815
rect -807 -1849 -773 -1825
rect -807 -1893 -773 -1887
rect -807 -1921 -773 -1893
rect -807 -1961 -773 -1959
rect -807 -1993 -773 -1961
rect -807 -2063 -773 -2031
rect -807 -2065 -773 -2063
rect -807 -2131 -773 -2103
rect -807 -2137 -773 -2131
rect -807 -2199 -773 -2175
rect -807 -2209 -773 -2199
rect -807 -2267 -773 -2247
rect -807 -2281 -773 -2267
rect -807 -2335 -773 -2319
rect -807 -2353 -773 -2335
rect -807 -2403 -773 -2391
rect -807 -2425 -773 -2403
rect -807 -2471 -773 -2463
rect -807 -2497 -773 -2471
rect -807 -2539 -773 -2535
rect -807 -2569 -773 -2539
rect -649 -1485 -615 -1455
rect -649 -1489 -615 -1485
rect -649 -1553 -615 -1527
rect -649 -1561 -615 -1553
rect -649 -1621 -615 -1599
rect -649 -1633 -615 -1621
rect -649 -1689 -615 -1671
rect -649 -1705 -615 -1689
rect -649 -1757 -615 -1743
rect -649 -1777 -615 -1757
rect -649 -1825 -615 -1815
rect -649 -1849 -615 -1825
rect -649 -1893 -615 -1887
rect -649 -1921 -615 -1893
rect -649 -1961 -615 -1959
rect -649 -1993 -615 -1961
rect -649 -2063 -615 -2031
rect -649 -2065 -615 -2063
rect -649 -2131 -615 -2103
rect -649 -2137 -615 -2131
rect -649 -2199 -615 -2175
rect -649 -2209 -615 -2199
rect -649 -2267 -615 -2247
rect -649 -2281 -615 -2267
rect -649 -2335 -615 -2319
rect -649 -2353 -615 -2335
rect -649 -2403 -615 -2391
rect -649 -2425 -615 -2403
rect -649 -2471 -615 -2463
rect -649 -2497 -615 -2471
rect -649 -2539 -615 -2535
rect -649 -2569 -615 -2539
rect -491 -1485 -457 -1455
rect -491 -1489 -457 -1485
rect -491 -1553 -457 -1527
rect -491 -1561 -457 -1553
rect -491 -1621 -457 -1599
rect -491 -1633 -457 -1621
rect -491 -1689 -457 -1671
rect -491 -1705 -457 -1689
rect -491 -1757 -457 -1743
rect -491 -1777 -457 -1757
rect -491 -1825 -457 -1815
rect -491 -1849 -457 -1825
rect -491 -1893 -457 -1887
rect -491 -1921 -457 -1893
rect -491 -1961 -457 -1959
rect -491 -1993 -457 -1961
rect -491 -2063 -457 -2031
rect -491 -2065 -457 -2063
rect -491 -2131 -457 -2103
rect -491 -2137 -457 -2131
rect -491 -2199 -457 -2175
rect -491 -2209 -457 -2199
rect -491 -2267 -457 -2247
rect -491 -2281 -457 -2267
rect -491 -2335 -457 -2319
rect -491 -2353 -457 -2335
rect -491 -2403 -457 -2391
rect -491 -2425 -457 -2403
rect -491 -2471 -457 -2463
rect -491 -2497 -457 -2471
rect -491 -2539 -457 -2535
rect -491 -2569 -457 -2539
rect -333 -1485 -299 -1455
rect -333 -1489 -299 -1485
rect -333 -1553 -299 -1527
rect -333 -1561 -299 -1553
rect -333 -1621 -299 -1599
rect -333 -1633 -299 -1621
rect -333 -1689 -299 -1671
rect -333 -1705 -299 -1689
rect -333 -1757 -299 -1743
rect -333 -1777 -299 -1757
rect -333 -1825 -299 -1815
rect -333 -1849 -299 -1825
rect -333 -1893 -299 -1887
rect -333 -1921 -299 -1893
rect -333 -1961 -299 -1959
rect -333 -1993 -299 -1961
rect -333 -2063 -299 -2031
rect -333 -2065 -299 -2063
rect -333 -2131 -299 -2103
rect -333 -2137 -299 -2131
rect -333 -2199 -299 -2175
rect -333 -2209 -299 -2199
rect -333 -2267 -299 -2247
rect -333 -2281 -299 -2267
rect -333 -2335 -299 -2319
rect -333 -2353 -299 -2335
rect -333 -2403 -299 -2391
rect -333 -2425 -299 -2403
rect -333 -2471 -299 -2463
rect -333 -2497 -299 -2471
rect -333 -2539 -299 -2535
rect -333 -2569 -299 -2539
rect -175 -1485 -141 -1455
rect -175 -1489 -141 -1485
rect -175 -1553 -141 -1527
rect -175 -1561 -141 -1553
rect -175 -1621 -141 -1599
rect -175 -1633 -141 -1621
rect -175 -1689 -141 -1671
rect -175 -1705 -141 -1689
rect -175 -1757 -141 -1743
rect -175 -1777 -141 -1757
rect -175 -1825 -141 -1815
rect -175 -1849 -141 -1825
rect -175 -1893 -141 -1887
rect -175 -1921 -141 -1893
rect -175 -1961 -141 -1959
rect -175 -1993 -141 -1961
rect -175 -2063 -141 -2031
rect -175 -2065 -141 -2063
rect -175 -2131 -141 -2103
rect -175 -2137 -141 -2131
rect -175 -2199 -141 -2175
rect -175 -2209 -141 -2199
rect -175 -2267 -141 -2247
rect -175 -2281 -141 -2267
rect -175 -2335 -141 -2319
rect -175 -2353 -141 -2335
rect -175 -2403 -141 -2391
rect -175 -2425 -141 -2403
rect -175 -2471 -141 -2463
rect -175 -2497 -141 -2471
rect -175 -2539 -141 -2535
rect -175 -2569 -141 -2539
rect -17 -1485 17 -1455
rect -17 -1489 17 -1485
rect -17 -1553 17 -1527
rect -17 -1561 17 -1553
rect -17 -1621 17 -1599
rect -17 -1633 17 -1621
rect -17 -1689 17 -1671
rect -17 -1705 17 -1689
rect -17 -1757 17 -1743
rect -17 -1777 17 -1757
rect -17 -1825 17 -1815
rect -17 -1849 17 -1825
rect -17 -1893 17 -1887
rect -17 -1921 17 -1893
rect -17 -1961 17 -1959
rect -17 -1993 17 -1961
rect -17 -2063 17 -2031
rect -17 -2065 17 -2063
rect -17 -2131 17 -2103
rect -17 -2137 17 -2131
rect -17 -2199 17 -2175
rect -17 -2209 17 -2199
rect -17 -2267 17 -2247
rect -17 -2281 17 -2267
rect -17 -2335 17 -2319
rect -17 -2353 17 -2335
rect -17 -2403 17 -2391
rect -17 -2425 17 -2403
rect -17 -2471 17 -2463
rect -17 -2497 17 -2471
rect -17 -2539 17 -2535
rect -17 -2569 17 -2539
rect 141 -1485 175 -1455
rect 141 -1489 175 -1485
rect 141 -1553 175 -1527
rect 141 -1561 175 -1553
rect 141 -1621 175 -1599
rect 141 -1633 175 -1621
rect 141 -1689 175 -1671
rect 141 -1705 175 -1689
rect 141 -1757 175 -1743
rect 141 -1777 175 -1757
rect 141 -1825 175 -1815
rect 141 -1849 175 -1825
rect 141 -1893 175 -1887
rect 141 -1921 175 -1893
rect 141 -1961 175 -1959
rect 141 -1993 175 -1961
rect 141 -2063 175 -2031
rect 141 -2065 175 -2063
rect 141 -2131 175 -2103
rect 141 -2137 175 -2131
rect 141 -2199 175 -2175
rect 141 -2209 175 -2199
rect 141 -2267 175 -2247
rect 141 -2281 175 -2267
rect 141 -2335 175 -2319
rect 141 -2353 175 -2335
rect 141 -2403 175 -2391
rect 141 -2425 175 -2403
rect 141 -2471 175 -2463
rect 141 -2497 175 -2471
rect 141 -2539 175 -2535
rect 141 -2569 175 -2539
rect 299 -1485 333 -1455
rect 299 -1489 333 -1485
rect 299 -1553 333 -1527
rect 299 -1561 333 -1553
rect 299 -1621 333 -1599
rect 299 -1633 333 -1621
rect 299 -1689 333 -1671
rect 299 -1705 333 -1689
rect 299 -1757 333 -1743
rect 299 -1777 333 -1757
rect 299 -1825 333 -1815
rect 299 -1849 333 -1825
rect 299 -1893 333 -1887
rect 299 -1921 333 -1893
rect 299 -1961 333 -1959
rect 299 -1993 333 -1961
rect 299 -2063 333 -2031
rect 299 -2065 333 -2063
rect 299 -2131 333 -2103
rect 299 -2137 333 -2131
rect 299 -2199 333 -2175
rect 299 -2209 333 -2199
rect 299 -2267 333 -2247
rect 299 -2281 333 -2267
rect 299 -2335 333 -2319
rect 299 -2353 333 -2335
rect 299 -2403 333 -2391
rect 299 -2425 333 -2403
rect 299 -2471 333 -2463
rect 299 -2497 333 -2471
rect 299 -2539 333 -2535
rect 299 -2569 333 -2539
rect 457 -1485 491 -1455
rect 457 -1489 491 -1485
rect 457 -1553 491 -1527
rect 457 -1561 491 -1553
rect 457 -1621 491 -1599
rect 457 -1633 491 -1621
rect 457 -1689 491 -1671
rect 457 -1705 491 -1689
rect 457 -1757 491 -1743
rect 457 -1777 491 -1757
rect 457 -1825 491 -1815
rect 457 -1849 491 -1825
rect 457 -1893 491 -1887
rect 457 -1921 491 -1893
rect 457 -1961 491 -1959
rect 457 -1993 491 -1961
rect 457 -2063 491 -2031
rect 457 -2065 491 -2063
rect 457 -2131 491 -2103
rect 457 -2137 491 -2131
rect 457 -2199 491 -2175
rect 457 -2209 491 -2199
rect 457 -2267 491 -2247
rect 457 -2281 491 -2267
rect 457 -2335 491 -2319
rect 457 -2353 491 -2335
rect 457 -2403 491 -2391
rect 457 -2425 491 -2403
rect 457 -2471 491 -2463
rect 457 -2497 491 -2471
rect 457 -2539 491 -2535
rect 457 -2569 491 -2539
rect 615 -1485 649 -1455
rect 615 -1489 649 -1485
rect 615 -1553 649 -1527
rect 615 -1561 649 -1553
rect 615 -1621 649 -1599
rect 615 -1633 649 -1621
rect 615 -1689 649 -1671
rect 615 -1705 649 -1689
rect 615 -1757 649 -1743
rect 615 -1777 649 -1757
rect 615 -1825 649 -1815
rect 615 -1849 649 -1825
rect 615 -1893 649 -1887
rect 615 -1921 649 -1893
rect 615 -1961 649 -1959
rect 615 -1993 649 -1961
rect 615 -2063 649 -2031
rect 615 -2065 649 -2063
rect 615 -2131 649 -2103
rect 615 -2137 649 -2131
rect 615 -2199 649 -2175
rect 615 -2209 649 -2199
rect 615 -2267 649 -2247
rect 615 -2281 649 -2267
rect 615 -2335 649 -2319
rect 615 -2353 649 -2335
rect 615 -2403 649 -2391
rect 615 -2425 649 -2403
rect 615 -2471 649 -2463
rect 615 -2497 649 -2471
rect 615 -2539 649 -2535
rect 615 -2569 649 -2539
rect 773 -1485 807 -1455
rect 773 -1489 807 -1485
rect 773 -1553 807 -1527
rect 773 -1561 807 -1553
rect 773 -1621 807 -1599
rect 773 -1633 807 -1621
rect 773 -1689 807 -1671
rect 773 -1705 807 -1689
rect 773 -1757 807 -1743
rect 773 -1777 807 -1757
rect 773 -1825 807 -1815
rect 773 -1849 807 -1825
rect 773 -1893 807 -1887
rect 773 -1921 807 -1893
rect 773 -1961 807 -1959
rect 773 -1993 807 -1961
rect 773 -2063 807 -2031
rect 773 -2065 807 -2063
rect 773 -2131 807 -2103
rect 773 -2137 807 -2131
rect 773 -2199 807 -2175
rect 773 -2209 807 -2199
rect 773 -2267 807 -2247
rect 773 -2281 807 -2267
rect 773 -2335 807 -2319
rect 773 -2353 807 -2335
rect 773 -2403 807 -2391
rect 773 -2425 807 -2403
rect 773 -2471 807 -2463
rect 773 -2497 807 -2471
rect 773 -2539 807 -2535
rect 773 -2569 807 -2539
rect 931 -1485 965 -1455
rect 931 -1489 965 -1485
rect 931 -1553 965 -1527
rect 931 -1561 965 -1553
rect 931 -1621 965 -1599
rect 931 -1633 965 -1621
rect 931 -1689 965 -1671
rect 931 -1705 965 -1689
rect 931 -1757 965 -1743
rect 931 -1777 965 -1757
rect 931 -1825 965 -1815
rect 931 -1849 965 -1825
rect 931 -1893 965 -1887
rect 931 -1921 965 -1893
rect 931 -1961 965 -1959
rect 931 -1993 965 -1961
rect 931 -2063 965 -2031
rect 931 -2065 965 -2063
rect 931 -2131 965 -2103
rect 931 -2137 965 -2131
rect 931 -2199 965 -2175
rect 931 -2209 965 -2199
rect 931 -2267 965 -2247
rect 931 -2281 965 -2267
rect 931 -2335 965 -2319
rect 931 -2353 965 -2335
rect 931 -2403 965 -2391
rect 931 -2425 965 -2403
rect 931 -2471 965 -2463
rect 931 -2497 965 -2471
rect 931 -2539 965 -2535
rect 931 -2569 965 -2539
rect 1089 -1485 1123 -1455
rect 1089 -1489 1123 -1485
rect 1089 -1553 1123 -1527
rect 1089 -1561 1123 -1553
rect 1089 -1621 1123 -1599
rect 1089 -1633 1123 -1621
rect 1089 -1689 1123 -1671
rect 1089 -1705 1123 -1689
rect 1089 -1757 1123 -1743
rect 1089 -1777 1123 -1757
rect 1089 -1825 1123 -1815
rect 1089 -1849 1123 -1825
rect 1089 -1893 1123 -1887
rect 1089 -1921 1123 -1893
rect 1089 -1961 1123 -1959
rect 1089 -1993 1123 -1961
rect 1089 -2063 1123 -2031
rect 1089 -2065 1123 -2063
rect 1089 -2131 1123 -2103
rect 1089 -2137 1123 -2131
rect 1089 -2199 1123 -2175
rect 1089 -2209 1123 -2199
rect 1089 -2267 1123 -2247
rect 1089 -2281 1123 -2267
rect 1089 -2335 1123 -2319
rect 1089 -2353 1123 -2335
rect 1089 -2403 1123 -2391
rect 1089 -2425 1123 -2403
rect 1089 -2471 1123 -2463
rect 1089 -2497 1123 -2471
rect 1089 -2539 1123 -2535
rect 1089 -2569 1123 -2539
rect -1044 -2693 -1010 -2659
rect -886 -2693 -852 -2659
rect -728 -2693 -694 -2659
rect -570 -2693 -536 -2659
rect -412 -2693 -378 -2659
rect -254 -2693 -220 -2659
rect -96 -2693 -62 -2659
rect 62 -2693 96 -2659
rect 220 -2693 254 -2659
rect 378 -2693 412 -2659
rect 536 -2693 570 -2659
rect 694 -2693 728 -2659
rect 852 -2693 886 -2659
rect 1010 -2693 1044 -2659
<< metal1 >>
rect -1129 2640 -1083 2683
rect -1129 2606 -1123 2640
rect -1089 2606 -1083 2640
rect -1129 2568 -1083 2606
rect -1129 2534 -1123 2568
rect -1089 2534 -1083 2568
rect -1129 2496 -1083 2534
rect -1129 2462 -1123 2496
rect -1089 2462 -1083 2496
rect -1129 2424 -1083 2462
rect -1129 2390 -1123 2424
rect -1089 2390 -1083 2424
rect -1129 2352 -1083 2390
rect -1129 2318 -1123 2352
rect -1089 2318 -1083 2352
rect -1129 2280 -1083 2318
rect -1129 2246 -1123 2280
rect -1089 2246 -1083 2280
rect -1129 2208 -1083 2246
rect -1129 2174 -1123 2208
rect -1089 2174 -1083 2208
rect -1129 2136 -1083 2174
rect -1129 2102 -1123 2136
rect -1089 2102 -1083 2136
rect -1129 2064 -1083 2102
rect -1129 2030 -1123 2064
rect -1089 2030 -1083 2064
rect -1129 1992 -1083 2030
rect -1129 1958 -1123 1992
rect -1089 1958 -1083 1992
rect -1129 1920 -1083 1958
rect -1129 1886 -1123 1920
rect -1089 1886 -1083 1920
rect -1129 1848 -1083 1886
rect -1129 1814 -1123 1848
rect -1089 1814 -1083 1848
rect -1129 1776 -1083 1814
rect -1129 1742 -1123 1776
rect -1089 1742 -1083 1776
rect -1129 1704 -1083 1742
rect -1129 1670 -1123 1704
rect -1089 1670 -1083 1704
rect -1129 1632 -1083 1670
rect -1129 1598 -1123 1632
rect -1089 1598 -1083 1632
rect -1129 1560 -1083 1598
rect -1129 1526 -1123 1560
rect -1089 1526 -1083 1560
rect -1129 1483 -1083 1526
rect -971 2640 -925 2683
rect -971 2606 -965 2640
rect -931 2606 -925 2640
rect -971 2568 -925 2606
rect -971 2534 -965 2568
rect -931 2534 -925 2568
rect -971 2496 -925 2534
rect -971 2462 -965 2496
rect -931 2462 -925 2496
rect -971 2424 -925 2462
rect -971 2390 -965 2424
rect -931 2390 -925 2424
rect -971 2352 -925 2390
rect -971 2318 -965 2352
rect -931 2318 -925 2352
rect -971 2280 -925 2318
rect -971 2246 -965 2280
rect -931 2246 -925 2280
rect -971 2208 -925 2246
rect -971 2174 -965 2208
rect -931 2174 -925 2208
rect -971 2136 -925 2174
rect -971 2102 -965 2136
rect -931 2102 -925 2136
rect -971 2064 -925 2102
rect -971 2030 -965 2064
rect -931 2030 -925 2064
rect -971 1992 -925 2030
rect -971 1958 -965 1992
rect -931 1958 -925 1992
rect -971 1920 -925 1958
rect -971 1886 -965 1920
rect -931 1886 -925 1920
rect -971 1848 -925 1886
rect -971 1814 -965 1848
rect -931 1814 -925 1848
rect -971 1776 -925 1814
rect -971 1742 -965 1776
rect -931 1742 -925 1776
rect -971 1704 -925 1742
rect -971 1670 -965 1704
rect -931 1670 -925 1704
rect -971 1632 -925 1670
rect -971 1598 -965 1632
rect -931 1598 -925 1632
rect -971 1560 -925 1598
rect -971 1526 -965 1560
rect -931 1526 -925 1560
rect -971 1483 -925 1526
rect -813 2640 -767 2683
rect -813 2606 -807 2640
rect -773 2606 -767 2640
rect -813 2568 -767 2606
rect -813 2534 -807 2568
rect -773 2534 -767 2568
rect -813 2496 -767 2534
rect -813 2462 -807 2496
rect -773 2462 -767 2496
rect -813 2424 -767 2462
rect -813 2390 -807 2424
rect -773 2390 -767 2424
rect -813 2352 -767 2390
rect -813 2318 -807 2352
rect -773 2318 -767 2352
rect -813 2280 -767 2318
rect -813 2246 -807 2280
rect -773 2246 -767 2280
rect -813 2208 -767 2246
rect -813 2174 -807 2208
rect -773 2174 -767 2208
rect -813 2136 -767 2174
rect -813 2102 -807 2136
rect -773 2102 -767 2136
rect -813 2064 -767 2102
rect -813 2030 -807 2064
rect -773 2030 -767 2064
rect -813 1992 -767 2030
rect -813 1958 -807 1992
rect -773 1958 -767 1992
rect -813 1920 -767 1958
rect -813 1886 -807 1920
rect -773 1886 -767 1920
rect -813 1848 -767 1886
rect -813 1814 -807 1848
rect -773 1814 -767 1848
rect -813 1776 -767 1814
rect -813 1742 -807 1776
rect -773 1742 -767 1776
rect -813 1704 -767 1742
rect -813 1670 -807 1704
rect -773 1670 -767 1704
rect -813 1632 -767 1670
rect -813 1598 -807 1632
rect -773 1598 -767 1632
rect -813 1560 -767 1598
rect -813 1526 -807 1560
rect -773 1526 -767 1560
rect -813 1483 -767 1526
rect -655 2640 -609 2683
rect -655 2606 -649 2640
rect -615 2606 -609 2640
rect -655 2568 -609 2606
rect -655 2534 -649 2568
rect -615 2534 -609 2568
rect -655 2496 -609 2534
rect -655 2462 -649 2496
rect -615 2462 -609 2496
rect -655 2424 -609 2462
rect -655 2390 -649 2424
rect -615 2390 -609 2424
rect -655 2352 -609 2390
rect -655 2318 -649 2352
rect -615 2318 -609 2352
rect -655 2280 -609 2318
rect -655 2246 -649 2280
rect -615 2246 -609 2280
rect -655 2208 -609 2246
rect -655 2174 -649 2208
rect -615 2174 -609 2208
rect -655 2136 -609 2174
rect -655 2102 -649 2136
rect -615 2102 -609 2136
rect -655 2064 -609 2102
rect -655 2030 -649 2064
rect -615 2030 -609 2064
rect -655 1992 -609 2030
rect -655 1958 -649 1992
rect -615 1958 -609 1992
rect -655 1920 -609 1958
rect -655 1886 -649 1920
rect -615 1886 -609 1920
rect -655 1848 -609 1886
rect -655 1814 -649 1848
rect -615 1814 -609 1848
rect -655 1776 -609 1814
rect -655 1742 -649 1776
rect -615 1742 -609 1776
rect -655 1704 -609 1742
rect -655 1670 -649 1704
rect -615 1670 -609 1704
rect -655 1632 -609 1670
rect -655 1598 -649 1632
rect -615 1598 -609 1632
rect -655 1560 -609 1598
rect -655 1526 -649 1560
rect -615 1526 -609 1560
rect -655 1483 -609 1526
rect -497 2640 -451 2683
rect -497 2606 -491 2640
rect -457 2606 -451 2640
rect -497 2568 -451 2606
rect -497 2534 -491 2568
rect -457 2534 -451 2568
rect -497 2496 -451 2534
rect -497 2462 -491 2496
rect -457 2462 -451 2496
rect -497 2424 -451 2462
rect -497 2390 -491 2424
rect -457 2390 -451 2424
rect -497 2352 -451 2390
rect -497 2318 -491 2352
rect -457 2318 -451 2352
rect -497 2280 -451 2318
rect -497 2246 -491 2280
rect -457 2246 -451 2280
rect -497 2208 -451 2246
rect -497 2174 -491 2208
rect -457 2174 -451 2208
rect -497 2136 -451 2174
rect -497 2102 -491 2136
rect -457 2102 -451 2136
rect -497 2064 -451 2102
rect -497 2030 -491 2064
rect -457 2030 -451 2064
rect -497 1992 -451 2030
rect -497 1958 -491 1992
rect -457 1958 -451 1992
rect -497 1920 -451 1958
rect -497 1886 -491 1920
rect -457 1886 -451 1920
rect -497 1848 -451 1886
rect -497 1814 -491 1848
rect -457 1814 -451 1848
rect -497 1776 -451 1814
rect -497 1742 -491 1776
rect -457 1742 -451 1776
rect -497 1704 -451 1742
rect -497 1670 -491 1704
rect -457 1670 -451 1704
rect -497 1632 -451 1670
rect -497 1598 -491 1632
rect -457 1598 -451 1632
rect -497 1560 -451 1598
rect -497 1526 -491 1560
rect -457 1526 -451 1560
rect -497 1483 -451 1526
rect -339 2640 -293 2683
rect -339 2606 -333 2640
rect -299 2606 -293 2640
rect -339 2568 -293 2606
rect -339 2534 -333 2568
rect -299 2534 -293 2568
rect -339 2496 -293 2534
rect -339 2462 -333 2496
rect -299 2462 -293 2496
rect -339 2424 -293 2462
rect -339 2390 -333 2424
rect -299 2390 -293 2424
rect -339 2352 -293 2390
rect -339 2318 -333 2352
rect -299 2318 -293 2352
rect -339 2280 -293 2318
rect -339 2246 -333 2280
rect -299 2246 -293 2280
rect -339 2208 -293 2246
rect -339 2174 -333 2208
rect -299 2174 -293 2208
rect -339 2136 -293 2174
rect -339 2102 -333 2136
rect -299 2102 -293 2136
rect -339 2064 -293 2102
rect -339 2030 -333 2064
rect -299 2030 -293 2064
rect -339 1992 -293 2030
rect -339 1958 -333 1992
rect -299 1958 -293 1992
rect -339 1920 -293 1958
rect -339 1886 -333 1920
rect -299 1886 -293 1920
rect -339 1848 -293 1886
rect -339 1814 -333 1848
rect -299 1814 -293 1848
rect -339 1776 -293 1814
rect -339 1742 -333 1776
rect -299 1742 -293 1776
rect -339 1704 -293 1742
rect -339 1670 -333 1704
rect -299 1670 -293 1704
rect -339 1632 -293 1670
rect -339 1598 -333 1632
rect -299 1598 -293 1632
rect -339 1560 -293 1598
rect -339 1526 -333 1560
rect -299 1526 -293 1560
rect -339 1483 -293 1526
rect -181 2640 -135 2683
rect -181 2606 -175 2640
rect -141 2606 -135 2640
rect -181 2568 -135 2606
rect -181 2534 -175 2568
rect -141 2534 -135 2568
rect -181 2496 -135 2534
rect -181 2462 -175 2496
rect -141 2462 -135 2496
rect -181 2424 -135 2462
rect -181 2390 -175 2424
rect -141 2390 -135 2424
rect -181 2352 -135 2390
rect -181 2318 -175 2352
rect -141 2318 -135 2352
rect -181 2280 -135 2318
rect -181 2246 -175 2280
rect -141 2246 -135 2280
rect -181 2208 -135 2246
rect -181 2174 -175 2208
rect -141 2174 -135 2208
rect -181 2136 -135 2174
rect -181 2102 -175 2136
rect -141 2102 -135 2136
rect -181 2064 -135 2102
rect -181 2030 -175 2064
rect -141 2030 -135 2064
rect -181 1992 -135 2030
rect -181 1958 -175 1992
rect -141 1958 -135 1992
rect -181 1920 -135 1958
rect -181 1886 -175 1920
rect -141 1886 -135 1920
rect -181 1848 -135 1886
rect -181 1814 -175 1848
rect -141 1814 -135 1848
rect -181 1776 -135 1814
rect -181 1742 -175 1776
rect -141 1742 -135 1776
rect -181 1704 -135 1742
rect -181 1670 -175 1704
rect -141 1670 -135 1704
rect -181 1632 -135 1670
rect -181 1598 -175 1632
rect -141 1598 -135 1632
rect -181 1560 -135 1598
rect -181 1526 -175 1560
rect -141 1526 -135 1560
rect -181 1483 -135 1526
rect -23 2640 23 2683
rect -23 2606 -17 2640
rect 17 2606 23 2640
rect -23 2568 23 2606
rect -23 2534 -17 2568
rect 17 2534 23 2568
rect -23 2496 23 2534
rect -23 2462 -17 2496
rect 17 2462 23 2496
rect -23 2424 23 2462
rect -23 2390 -17 2424
rect 17 2390 23 2424
rect -23 2352 23 2390
rect -23 2318 -17 2352
rect 17 2318 23 2352
rect -23 2280 23 2318
rect -23 2246 -17 2280
rect 17 2246 23 2280
rect -23 2208 23 2246
rect -23 2174 -17 2208
rect 17 2174 23 2208
rect -23 2136 23 2174
rect -23 2102 -17 2136
rect 17 2102 23 2136
rect -23 2064 23 2102
rect -23 2030 -17 2064
rect 17 2030 23 2064
rect -23 1992 23 2030
rect -23 1958 -17 1992
rect 17 1958 23 1992
rect -23 1920 23 1958
rect -23 1886 -17 1920
rect 17 1886 23 1920
rect -23 1848 23 1886
rect -23 1814 -17 1848
rect 17 1814 23 1848
rect -23 1776 23 1814
rect -23 1742 -17 1776
rect 17 1742 23 1776
rect -23 1704 23 1742
rect -23 1670 -17 1704
rect 17 1670 23 1704
rect -23 1632 23 1670
rect -23 1598 -17 1632
rect 17 1598 23 1632
rect -23 1560 23 1598
rect -23 1526 -17 1560
rect 17 1526 23 1560
rect -23 1483 23 1526
rect 135 2640 181 2683
rect 135 2606 141 2640
rect 175 2606 181 2640
rect 135 2568 181 2606
rect 135 2534 141 2568
rect 175 2534 181 2568
rect 135 2496 181 2534
rect 135 2462 141 2496
rect 175 2462 181 2496
rect 135 2424 181 2462
rect 135 2390 141 2424
rect 175 2390 181 2424
rect 135 2352 181 2390
rect 135 2318 141 2352
rect 175 2318 181 2352
rect 135 2280 181 2318
rect 135 2246 141 2280
rect 175 2246 181 2280
rect 135 2208 181 2246
rect 135 2174 141 2208
rect 175 2174 181 2208
rect 135 2136 181 2174
rect 135 2102 141 2136
rect 175 2102 181 2136
rect 135 2064 181 2102
rect 135 2030 141 2064
rect 175 2030 181 2064
rect 135 1992 181 2030
rect 135 1958 141 1992
rect 175 1958 181 1992
rect 135 1920 181 1958
rect 135 1886 141 1920
rect 175 1886 181 1920
rect 135 1848 181 1886
rect 135 1814 141 1848
rect 175 1814 181 1848
rect 135 1776 181 1814
rect 135 1742 141 1776
rect 175 1742 181 1776
rect 135 1704 181 1742
rect 135 1670 141 1704
rect 175 1670 181 1704
rect 135 1632 181 1670
rect 135 1598 141 1632
rect 175 1598 181 1632
rect 135 1560 181 1598
rect 135 1526 141 1560
rect 175 1526 181 1560
rect 135 1483 181 1526
rect 293 2640 339 2683
rect 293 2606 299 2640
rect 333 2606 339 2640
rect 293 2568 339 2606
rect 293 2534 299 2568
rect 333 2534 339 2568
rect 293 2496 339 2534
rect 293 2462 299 2496
rect 333 2462 339 2496
rect 293 2424 339 2462
rect 293 2390 299 2424
rect 333 2390 339 2424
rect 293 2352 339 2390
rect 293 2318 299 2352
rect 333 2318 339 2352
rect 293 2280 339 2318
rect 293 2246 299 2280
rect 333 2246 339 2280
rect 293 2208 339 2246
rect 293 2174 299 2208
rect 333 2174 339 2208
rect 293 2136 339 2174
rect 293 2102 299 2136
rect 333 2102 339 2136
rect 293 2064 339 2102
rect 293 2030 299 2064
rect 333 2030 339 2064
rect 293 1992 339 2030
rect 293 1958 299 1992
rect 333 1958 339 1992
rect 293 1920 339 1958
rect 293 1886 299 1920
rect 333 1886 339 1920
rect 293 1848 339 1886
rect 293 1814 299 1848
rect 333 1814 339 1848
rect 293 1776 339 1814
rect 293 1742 299 1776
rect 333 1742 339 1776
rect 293 1704 339 1742
rect 293 1670 299 1704
rect 333 1670 339 1704
rect 293 1632 339 1670
rect 293 1598 299 1632
rect 333 1598 339 1632
rect 293 1560 339 1598
rect 293 1526 299 1560
rect 333 1526 339 1560
rect 293 1483 339 1526
rect 451 2640 497 2683
rect 451 2606 457 2640
rect 491 2606 497 2640
rect 451 2568 497 2606
rect 451 2534 457 2568
rect 491 2534 497 2568
rect 451 2496 497 2534
rect 451 2462 457 2496
rect 491 2462 497 2496
rect 451 2424 497 2462
rect 451 2390 457 2424
rect 491 2390 497 2424
rect 451 2352 497 2390
rect 451 2318 457 2352
rect 491 2318 497 2352
rect 451 2280 497 2318
rect 451 2246 457 2280
rect 491 2246 497 2280
rect 451 2208 497 2246
rect 451 2174 457 2208
rect 491 2174 497 2208
rect 451 2136 497 2174
rect 451 2102 457 2136
rect 491 2102 497 2136
rect 451 2064 497 2102
rect 451 2030 457 2064
rect 491 2030 497 2064
rect 451 1992 497 2030
rect 451 1958 457 1992
rect 491 1958 497 1992
rect 451 1920 497 1958
rect 451 1886 457 1920
rect 491 1886 497 1920
rect 451 1848 497 1886
rect 451 1814 457 1848
rect 491 1814 497 1848
rect 451 1776 497 1814
rect 451 1742 457 1776
rect 491 1742 497 1776
rect 451 1704 497 1742
rect 451 1670 457 1704
rect 491 1670 497 1704
rect 451 1632 497 1670
rect 451 1598 457 1632
rect 491 1598 497 1632
rect 451 1560 497 1598
rect 451 1526 457 1560
rect 491 1526 497 1560
rect 451 1483 497 1526
rect 609 2640 655 2683
rect 609 2606 615 2640
rect 649 2606 655 2640
rect 609 2568 655 2606
rect 609 2534 615 2568
rect 649 2534 655 2568
rect 609 2496 655 2534
rect 609 2462 615 2496
rect 649 2462 655 2496
rect 609 2424 655 2462
rect 609 2390 615 2424
rect 649 2390 655 2424
rect 609 2352 655 2390
rect 609 2318 615 2352
rect 649 2318 655 2352
rect 609 2280 655 2318
rect 609 2246 615 2280
rect 649 2246 655 2280
rect 609 2208 655 2246
rect 609 2174 615 2208
rect 649 2174 655 2208
rect 609 2136 655 2174
rect 609 2102 615 2136
rect 649 2102 655 2136
rect 609 2064 655 2102
rect 609 2030 615 2064
rect 649 2030 655 2064
rect 609 1992 655 2030
rect 609 1958 615 1992
rect 649 1958 655 1992
rect 609 1920 655 1958
rect 609 1886 615 1920
rect 649 1886 655 1920
rect 609 1848 655 1886
rect 609 1814 615 1848
rect 649 1814 655 1848
rect 609 1776 655 1814
rect 609 1742 615 1776
rect 649 1742 655 1776
rect 609 1704 655 1742
rect 609 1670 615 1704
rect 649 1670 655 1704
rect 609 1632 655 1670
rect 609 1598 615 1632
rect 649 1598 655 1632
rect 609 1560 655 1598
rect 609 1526 615 1560
rect 649 1526 655 1560
rect 609 1483 655 1526
rect 767 2640 813 2683
rect 767 2606 773 2640
rect 807 2606 813 2640
rect 767 2568 813 2606
rect 767 2534 773 2568
rect 807 2534 813 2568
rect 767 2496 813 2534
rect 767 2462 773 2496
rect 807 2462 813 2496
rect 767 2424 813 2462
rect 767 2390 773 2424
rect 807 2390 813 2424
rect 767 2352 813 2390
rect 767 2318 773 2352
rect 807 2318 813 2352
rect 767 2280 813 2318
rect 767 2246 773 2280
rect 807 2246 813 2280
rect 767 2208 813 2246
rect 767 2174 773 2208
rect 807 2174 813 2208
rect 767 2136 813 2174
rect 767 2102 773 2136
rect 807 2102 813 2136
rect 767 2064 813 2102
rect 767 2030 773 2064
rect 807 2030 813 2064
rect 767 1992 813 2030
rect 767 1958 773 1992
rect 807 1958 813 1992
rect 767 1920 813 1958
rect 767 1886 773 1920
rect 807 1886 813 1920
rect 767 1848 813 1886
rect 767 1814 773 1848
rect 807 1814 813 1848
rect 767 1776 813 1814
rect 767 1742 773 1776
rect 807 1742 813 1776
rect 767 1704 813 1742
rect 767 1670 773 1704
rect 807 1670 813 1704
rect 767 1632 813 1670
rect 767 1598 773 1632
rect 807 1598 813 1632
rect 767 1560 813 1598
rect 767 1526 773 1560
rect 807 1526 813 1560
rect 767 1483 813 1526
rect 925 2640 971 2683
rect 925 2606 931 2640
rect 965 2606 971 2640
rect 925 2568 971 2606
rect 925 2534 931 2568
rect 965 2534 971 2568
rect 925 2496 971 2534
rect 925 2462 931 2496
rect 965 2462 971 2496
rect 925 2424 971 2462
rect 925 2390 931 2424
rect 965 2390 971 2424
rect 925 2352 971 2390
rect 925 2318 931 2352
rect 965 2318 971 2352
rect 925 2280 971 2318
rect 925 2246 931 2280
rect 965 2246 971 2280
rect 925 2208 971 2246
rect 925 2174 931 2208
rect 965 2174 971 2208
rect 925 2136 971 2174
rect 925 2102 931 2136
rect 965 2102 971 2136
rect 925 2064 971 2102
rect 925 2030 931 2064
rect 965 2030 971 2064
rect 925 1992 971 2030
rect 925 1958 931 1992
rect 965 1958 971 1992
rect 925 1920 971 1958
rect 925 1886 931 1920
rect 965 1886 971 1920
rect 925 1848 971 1886
rect 925 1814 931 1848
rect 965 1814 971 1848
rect 925 1776 971 1814
rect 925 1742 931 1776
rect 965 1742 971 1776
rect 925 1704 971 1742
rect 925 1670 931 1704
rect 965 1670 971 1704
rect 925 1632 971 1670
rect 925 1598 931 1632
rect 965 1598 971 1632
rect 925 1560 971 1598
rect 925 1526 931 1560
rect 965 1526 971 1560
rect 925 1483 971 1526
rect 1083 2640 1129 2683
rect 1083 2606 1089 2640
rect 1123 2606 1129 2640
rect 1083 2568 1129 2606
rect 1083 2534 1089 2568
rect 1123 2534 1129 2568
rect 1083 2496 1129 2534
rect 1083 2462 1089 2496
rect 1123 2462 1129 2496
rect 1083 2424 1129 2462
rect 1083 2390 1089 2424
rect 1123 2390 1129 2424
rect 1083 2352 1129 2390
rect 1083 2318 1089 2352
rect 1123 2318 1129 2352
rect 1083 2280 1129 2318
rect 1083 2246 1089 2280
rect 1123 2246 1129 2280
rect 1083 2208 1129 2246
rect 1083 2174 1089 2208
rect 1123 2174 1129 2208
rect 1083 2136 1129 2174
rect 1083 2102 1089 2136
rect 1123 2102 1129 2136
rect 1083 2064 1129 2102
rect 1083 2030 1089 2064
rect 1123 2030 1129 2064
rect 1083 1992 1129 2030
rect 1083 1958 1089 1992
rect 1123 1958 1129 1992
rect 1083 1920 1129 1958
rect 1083 1886 1089 1920
rect 1123 1886 1129 1920
rect 1083 1848 1129 1886
rect 1083 1814 1089 1848
rect 1123 1814 1129 1848
rect 1083 1776 1129 1814
rect 1083 1742 1089 1776
rect 1123 1742 1129 1776
rect 1083 1704 1129 1742
rect 1083 1670 1089 1704
rect 1123 1670 1129 1704
rect 1083 1632 1129 1670
rect 1083 1598 1089 1632
rect 1123 1598 1129 1632
rect 1083 1560 1129 1598
rect 1083 1526 1089 1560
rect 1123 1526 1129 1560
rect 1083 1483 1129 1526
rect -1073 1436 -981 1442
rect -1073 1402 -1044 1436
rect -1010 1402 -981 1436
rect -1073 1396 -981 1402
rect -915 1436 -823 1442
rect -915 1402 -886 1436
rect -852 1402 -823 1436
rect -915 1396 -823 1402
rect -757 1436 -665 1442
rect -757 1402 -728 1436
rect -694 1402 -665 1436
rect -757 1396 -665 1402
rect -599 1436 -507 1442
rect -599 1402 -570 1436
rect -536 1402 -507 1436
rect -599 1396 -507 1402
rect -441 1436 -349 1442
rect -441 1402 -412 1436
rect -378 1402 -349 1436
rect -441 1396 -349 1402
rect -283 1436 -191 1442
rect -283 1402 -254 1436
rect -220 1402 -191 1436
rect -283 1396 -191 1402
rect -125 1436 -33 1442
rect -125 1402 -96 1436
rect -62 1402 -33 1436
rect -125 1396 -33 1402
rect 33 1436 125 1442
rect 33 1402 62 1436
rect 96 1402 125 1436
rect 33 1396 125 1402
rect 191 1436 283 1442
rect 191 1402 220 1436
rect 254 1402 283 1436
rect 191 1396 283 1402
rect 349 1436 441 1442
rect 349 1402 378 1436
rect 412 1402 441 1436
rect 349 1396 441 1402
rect 507 1436 599 1442
rect 507 1402 536 1436
rect 570 1402 599 1436
rect 507 1396 599 1402
rect 665 1436 757 1442
rect 665 1402 694 1436
rect 728 1402 757 1436
rect 665 1396 757 1402
rect 823 1436 915 1442
rect 823 1402 852 1436
rect 886 1402 915 1436
rect 823 1396 915 1402
rect 981 1436 1073 1442
rect 981 1402 1010 1436
rect 1044 1402 1073 1436
rect 981 1396 1073 1402
rect -1129 1275 -1083 1318
rect -1129 1241 -1123 1275
rect -1089 1241 -1083 1275
rect -1129 1203 -1083 1241
rect -1129 1169 -1123 1203
rect -1089 1169 -1083 1203
rect -1129 1131 -1083 1169
rect -1129 1097 -1123 1131
rect -1089 1097 -1083 1131
rect -1129 1059 -1083 1097
rect -1129 1025 -1123 1059
rect -1089 1025 -1083 1059
rect -1129 987 -1083 1025
rect -1129 953 -1123 987
rect -1089 953 -1083 987
rect -1129 915 -1083 953
rect -1129 881 -1123 915
rect -1089 881 -1083 915
rect -1129 843 -1083 881
rect -1129 809 -1123 843
rect -1089 809 -1083 843
rect -1129 771 -1083 809
rect -1129 737 -1123 771
rect -1089 737 -1083 771
rect -1129 699 -1083 737
rect -1129 665 -1123 699
rect -1089 665 -1083 699
rect -1129 627 -1083 665
rect -1129 593 -1123 627
rect -1089 593 -1083 627
rect -1129 555 -1083 593
rect -1129 521 -1123 555
rect -1089 521 -1083 555
rect -1129 483 -1083 521
rect -1129 449 -1123 483
rect -1089 449 -1083 483
rect -1129 411 -1083 449
rect -1129 377 -1123 411
rect -1089 377 -1083 411
rect -1129 339 -1083 377
rect -1129 305 -1123 339
rect -1089 305 -1083 339
rect -1129 267 -1083 305
rect -1129 233 -1123 267
rect -1089 233 -1083 267
rect -1129 195 -1083 233
rect -1129 161 -1123 195
rect -1089 161 -1083 195
rect -1129 118 -1083 161
rect -971 1275 -925 1318
rect -971 1241 -965 1275
rect -931 1241 -925 1275
rect -971 1203 -925 1241
rect -971 1169 -965 1203
rect -931 1169 -925 1203
rect -971 1131 -925 1169
rect -971 1097 -965 1131
rect -931 1097 -925 1131
rect -971 1059 -925 1097
rect -971 1025 -965 1059
rect -931 1025 -925 1059
rect -971 987 -925 1025
rect -971 953 -965 987
rect -931 953 -925 987
rect -971 915 -925 953
rect -971 881 -965 915
rect -931 881 -925 915
rect -971 843 -925 881
rect -971 809 -965 843
rect -931 809 -925 843
rect -971 771 -925 809
rect -971 737 -965 771
rect -931 737 -925 771
rect -971 699 -925 737
rect -971 665 -965 699
rect -931 665 -925 699
rect -971 627 -925 665
rect -971 593 -965 627
rect -931 593 -925 627
rect -971 555 -925 593
rect -971 521 -965 555
rect -931 521 -925 555
rect -971 483 -925 521
rect -971 449 -965 483
rect -931 449 -925 483
rect -971 411 -925 449
rect -971 377 -965 411
rect -931 377 -925 411
rect -971 339 -925 377
rect -971 305 -965 339
rect -931 305 -925 339
rect -971 267 -925 305
rect -971 233 -965 267
rect -931 233 -925 267
rect -971 195 -925 233
rect -971 161 -965 195
rect -931 161 -925 195
rect -971 118 -925 161
rect -813 1275 -767 1318
rect -813 1241 -807 1275
rect -773 1241 -767 1275
rect -813 1203 -767 1241
rect -813 1169 -807 1203
rect -773 1169 -767 1203
rect -813 1131 -767 1169
rect -813 1097 -807 1131
rect -773 1097 -767 1131
rect -813 1059 -767 1097
rect -813 1025 -807 1059
rect -773 1025 -767 1059
rect -813 987 -767 1025
rect -813 953 -807 987
rect -773 953 -767 987
rect -813 915 -767 953
rect -813 881 -807 915
rect -773 881 -767 915
rect -813 843 -767 881
rect -813 809 -807 843
rect -773 809 -767 843
rect -813 771 -767 809
rect -813 737 -807 771
rect -773 737 -767 771
rect -813 699 -767 737
rect -813 665 -807 699
rect -773 665 -767 699
rect -813 627 -767 665
rect -813 593 -807 627
rect -773 593 -767 627
rect -813 555 -767 593
rect -813 521 -807 555
rect -773 521 -767 555
rect -813 483 -767 521
rect -813 449 -807 483
rect -773 449 -767 483
rect -813 411 -767 449
rect -813 377 -807 411
rect -773 377 -767 411
rect -813 339 -767 377
rect -813 305 -807 339
rect -773 305 -767 339
rect -813 267 -767 305
rect -813 233 -807 267
rect -773 233 -767 267
rect -813 195 -767 233
rect -813 161 -807 195
rect -773 161 -767 195
rect -813 118 -767 161
rect -655 1275 -609 1318
rect -655 1241 -649 1275
rect -615 1241 -609 1275
rect -655 1203 -609 1241
rect -655 1169 -649 1203
rect -615 1169 -609 1203
rect -655 1131 -609 1169
rect -655 1097 -649 1131
rect -615 1097 -609 1131
rect -655 1059 -609 1097
rect -655 1025 -649 1059
rect -615 1025 -609 1059
rect -655 987 -609 1025
rect -655 953 -649 987
rect -615 953 -609 987
rect -655 915 -609 953
rect -655 881 -649 915
rect -615 881 -609 915
rect -655 843 -609 881
rect -655 809 -649 843
rect -615 809 -609 843
rect -655 771 -609 809
rect -655 737 -649 771
rect -615 737 -609 771
rect -655 699 -609 737
rect -655 665 -649 699
rect -615 665 -609 699
rect -655 627 -609 665
rect -655 593 -649 627
rect -615 593 -609 627
rect -655 555 -609 593
rect -655 521 -649 555
rect -615 521 -609 555
rect -655 483 -609 521
rect -655 449 -649 483
rect -615 449 -609 483
rect -655 411 -609 449
rect -655 377 -649 411
rect -615 377 -609 411
rect -655 339 -609 377
rect -655 305 -649 339
rect -615 305 -609 339
rect -655 267 -609 305
rect -655 233 -649 267
rect -615 233 -609 267
rect -655 195 -609 233
rect -655 161 -649 195
rect -615 161 -609 195
rect -655 118 -609 161
rect -497 1275 -451 1318
rect -497 1241 -491 1275
rect -457 1241 -451 1275
rect -497 1203 -451 1241
rect -497 1169 -491 1203
rect -457 1169 -451 1203
rect -497 1131 -451 1169
rect -497 1097 -491 1131
rect -457 1097 -451 1131
rect -497 1059 -451 1097
rect -497 1025 -491 1059
rect -457 1025 -451 1059
rect -497 987 -451 1025
rect -497 953 -491 987
rect -457 953 -451 987
rect -497 915 -451 953
rect -497 881 -491 915
rect -457 881 -451 915
rect -497 843 -451 881
rect -497 809 -491 843
rect -457 809 -451 843
rect -497 771 -451 809
rect -497 737 -491 771
rect -457 737 -451 771
rect -497 699 -451 737
rect -497 665 -491 699
rect -457 665 -451 699
rect -497 627 -451 665
rect -497 593 -491 627
rect -457 593 -451 627
rect -497 555 -451 593
rect -497 521 -491 555
rect -457 521 -451 555
rect -497 483 -451 521
rect -497 449 -491 483
rect -457 449 -451 483
rect -497 411 -451 449
rect -497 377 -491 411
rect -457 377 -451 411
rect -497 339 -451 377
rect -497 305 -491 339
rect -457 305 -451 339
rect -497 267 -451 305
rect -497 233 -491 267
rect -457 233 -451 267
rect -497 195 -451 233
rect -497 161 -491 195
rect -457 161 -451 195
rect -497 118 -451 161
rect -339 1275 -293 1318
rect -339 1241 -333 1275
rect -299 1241 -293 1275
rect -339 1203 -293 1241
rect -339 1169 -333 1203
rect -299 1169 -293 1203
rect -339 1131 -293 1169
rect -339 1097 -333 1131
rect -299 1097 -293 1131
rect -339 1059 -293 1097
rect -339 1025 -333 1059
rect -299 1025 -293 1059
rect -339 987 -293 1025
rect -339 953 -333 987
rect -299 953 -293 987
rect -339 915 -293 953
rect -339 881 -333 915
rect -299 881 -293 915
rect -339 843 -293 881
rect -339 809 -333 843
rect -299 809 -293 843
rect -339 771 -293 809
rect -339 737 -333 771
rect -299 737 -293 771
rect -339 699 -293 737
rect -339 665 -333 699
rect -299 665 -293 699
rect -339 627 -293 665
rect -339 593 -333 627
rect -299 593 -293 627
rect -339 555 -293 593
rect -339 521 -333 555
rect -299 521 -293 555
rect -339 483 -293 521
rect -339 449 -333 483
rect -299 449 -293 483
rect -339 411 -293 449
rect -339 377 -333 411
rect -299 377 -293 411
rect -339 339 -293 377
rect -339 305 -333 339
rect -299 305 -293 339
rect -339 267 -293 305
rect -339 233 -333 267
rect -299 233 -293 267
rect -339 195 -293 233
rect -339 161 -333 195
rect -299 161 -293 195
rect -339 118 -293 161
rect -181 1275 -135 1318
rect -181 1241 -175 1275
rect -141 1241 -135 1275
rect -181 1203 -135 1241
rect -181 1169 -175 1203
rect -141 1169 -135 1203
rect -181 1131 -135 1169
rect -181 1097 -175 1131
rect -141 1097 -135 1131
rect -181 1059 -135 1097
rect -181 1025 -175 1059
rect -141 1025 -135 1059
rect -181 987 -135 1025
rect -181 953 -175 987
rect -141 953 -135 987
rect -181 915 -135 953
rect -181 881 -175 915
rect -141 881 -135 915
rect -181 843 -135 881
rect -181 809 -175 843
rect -141 809 -135 843
rect -181 771 -135 809
rect -181 737 -175 771
rect -141 737 -135 771
rect -181 699 -135 737
rect -181 665 -175 699
rect -141 665 -135 699
rect -181 627 -135 665
rect -181 593 -175 627
rect -141 593 -135 627
rect -181 555 -135 593
rect -181 521 -175 555
rect -141 521 -135 555
rect -181 483 -135 521
rect -181 449 -175 483
rect -141 449 -135 483
rect -181 411 -135 449
rect -181 377 -175 411
rect -141 377 -135 411
rect -181 339 -135 377
rect -181 305 -175 339
rect -141 305 -135 339
rect -181 267 -135 305
rect -181 233 -175 267
rect -141 233 -135 267
rect -181 195 -135 233
rect -181 161 -175 195
rect -141 161 -135 195
rect -181 118 -135 161
rect -23 1275 23 1318
rect -23 1241 -17 1275
rect 17 1241 23 1275
rect -23 1203 23 1241
rect -23 1169 -17 1203
rect 17 1169 23 1203
rect -23 1131 23 1169
rect -23 1097 -17 1131
rect 17 1097 23 1131
rect -23 1059 23 1097
rect -23 1025 -17 1059
rect 17 1025 23 1059
rect -23 987 23 1025
rect -23 953 -17 987
rect 17 953 23 987
rect -23 915 23 953
rect -23 881 -17 915
rect 17 881 23 915
rect -23 843 23 881
rect -23 809 -17 843
rect 17 809 23 843
rect -23 771 23 809
rect -23 737 -17 771
rect 17 737 23 771
rect -23 699 23 737
rect -23 665 -17 699
rect 17 665 23 699
rect -23 627 23 665
rect -23 593 -17 627
rect 17 593 23 627
rect -23 555 23 593
rect -23 521 -17 555
rect 17 521 23 555
rect -23 483 23 521
rect -23 449 -17 483
rect 17 449 23 483
rect -23 411 23 449
rect -23 377 -17 411
rect 17 377 23 411
rect -23 339 23 377
rect -23 305 -17 339
rect 17 305 23 339
rect -23 267 23 305
rect -23 233 -17 267
rect 17 233 23 267
rect -23 195 23 233
rect -23 161 -17 195
rect 17 161 23 195
rect -23 118 23 161
rect 135 1275 181 1318
rect 135 1241 141 1275
rect 175 1241 181 1275
rect 135 1203 181 1241
rect 135 1169 141 1203
rect 175 1169 181 1203
rect 135 1131 181 1169
rect 135 1097 141 1131
rect 175 1097 181 1131
rect 135 1059 181 1097
rect 135 1025 141 1059
rect 175 1025 181 1059
rect 135 987 181 1025
rect 135 953 141 987
rect 175 953 181 987
rect 135 915 181 953
rect 135 881 141 915
rect 175 881 181 915
rect 135 843 181 881
rect 135 809 141 843
rect 175 809 181 843
rect 135 771 181 809
rect 135 737 141 771
rect 175 737 181 771
rect 135 699 181 737
rect 135 665 141 699
rect 175 665 181 699
rect 135 627 181 665
rect 135 593 141 627
rect 175 593 181 627
rect 135 555 181 593
rect 135 521 141 555
rect 175 521 181 555
rect 135 483 181 521
rect 135 449 141 483
rect 175 449 181 483
rect 135 411 181 449
rect 135 377 141 411
rect 175 377 181 411
rect 135 339 181 377
rect 135 305 141 339
rect 175 305 181 339
rect 135 267 181 305
rect 135 233 141 267
rect 175 233 181 267
rect 135 195 181 233
rect 135 161 141 195
rect 175 161 181 195
rect 135 118 181 161
rect 293 1275 339 1318
rect 293 1241 299 1275
rect 333 1241 339 1275
rect 293 1203 339 1241
rect 293 1169 299 1203
rect 333 1169 339 1203
rect 293 1131 339 1169
rect 293 1097 299 1131
rect 333 1097 339 1131
rect 293 1059 339 1097
rect 293 1025 299 1059
rect 333 1025 339 1059
rect 293 987 339 1025
rect 293 953 299 987
rect 333 953 339 987
rect 293 915 339 953
rect 293 881 299 915
rect 333 881 339 915
rect 293 843 339 881
rect 293 809 299 843
rect 333 809 339 843
rect 293 771 339 809
rect 293 737 299 771
rect 333 737 339 771
rect 293 699 339 737
rect 293 665 299 699
rect 333 665 339 699
rect 293 627 339 665
rect 293 593 299 627
rect 333 593 339 627
rect 293 555 339 593
rect 293 521 299 555
rect 333 521 339 555
rect 293 483 339 521
rect 293 449 299 483
rect 333 449 339 483
rect 293 411 339 449
rect 293 377 299 411
rect 333 377 339 411
rect 293 339 339 377
rect 293 305 299 339
rect 333 305 339 339
rect 293 267 339 305
rect 293 233 299 267
rect 333 233 339 267
rect 293 195 339 233
rect 293 161 299 195
rect 333 161 339 195
rect 293 118 339 161
rect 451 1275 497 1318
rect 451 1241 457 1275
rect 491 1241 497 1275
rect 451 1203 497 1241
rect 451 1169 457 1203
rect 491 1169 497 1203
rect 451 1131 497 1169
rect 451 1097 457 1131
rect 491 1097 497 1131
rect 451 1059 497 1097
rect 451 1025 457 1059
rect 491 1025 497 1059
rect 451 987 497 1025
rect 451 953 457 987
rect 491 953 497 987
rect 451 915 497 953
rect 451 881 457 915
rect 491 881 497 915
rect 451 843 497 881
rect 451 809 457 843
rect 491 809 497 843
rect 451 771 497 809
rect 451 737 457 771
rect 491 737 497 771
rect 451 699 497 737
rect 451 665 457 699
rect 491 665 497 699
rect 451 627 497 665
rect 451 593 457 627
rect 491 593 497 627
rect 451 555 497 593
rect 451 521 457 555
rect 491 521 497 555
rect 451 483 497 521
rect 451 449 457 483
rect 491 449 497 483
rect 451 411 497 449
rect 451 377 457 411
rect 491 377 497 411
rect 451 339 497 377
rect 451 305 457 339
rect 491 305 497 339
rect 451 267 497 305
rect 451 233 457 267
rect 491 233 497 267
rect 451 195 497 233
rect 451 161 457 195
rect 491 161 497 195
rect 451 118 497 161
rect 609 1275 655 1318
rect 609 1241 615 1275
rect 649 1241 655 1275
rect 609 1203 655 1241
rect 609 1169 615 1203
rect 649 1169 655 1203
rect 609 1131 655 1169
rect 609 1097 615 1131
rect 649 1097 655 1131
rect 609 1059 655 1097
rect 609 1025 615 1059
rect 649 1025 655 1059
rect 609 987 655 1025
rect 609 953 615 987
rect 649 953 655 987
rect 609 915 655 953
rect 609 881 615 915
rect 649 881 655 915
rect 609 843 655 881
rect 609 809 615 843
rect 649 809 655 843
rect 609 771 655 809
rect 609 737 615 771
rect 649 737 655 771
rect 609 699 655 737
rect 609 665 615 699
rect 649 665 655 699
rect 609 627 655 665
rect 609 593 615 627
rect 649 593 655 627
rect 609 555 655 593
rect 609 521 615 555
rect 649 521 655 555
rect 609 483 655 521
rect 609 449 615 483
rect 649 449 655 483
rect 609 411 655 449
rect 609 377 615 411
rect 649 377 655 411
rect 609 339 655 377
rect 609 305 615 339
rect 649 305 655 339
rect 609 267 655 305
rect 609 233 615 267
rect 649 233 655 267
rect 609 195 655 233
rect 609 161 615 195
rect 649 161 655 195
rect 609 118 655 161
rect 767 1275 813 1318
rect 767 1241 773 1275
rect 807 1241 813 1275
rect 767 1203 813 1241
rect 767 1169 773 1203
rect 807 1169 813 1203
rect 767 1131 813 1169
rect 767 1097 773 1131
rect 807 1097 813 1131
rect 767 1059 813 1097
rect 767 1025 773 1059
rect 807 1025 813 1059
rect 767 987 813 1025
rect 767 953 773 987
rect 807 953 813 987
rect 767 915 813 953
rect 767 881 773 915
rect 807 881 813 915
rect 767 843 813 881
rect 767 809 773 843
rect 807 809 813 843
rect 767 771 813 809
rect 767 737 773 771
rect 807 737 813 771
rect 767 699 813 737
rect 767 665 773 699
rect 807 665 813 699
rect 767 627 813 665
rect 767 593 773 627
rect 807 593 813 627
rect 767 555 813 593
rect 767 521 773 555
rect 807 521 813 555
rect 767 483 813 521
rect 767 449 773 483
rect 807 449 813 483
rect 767 411 813 449
rect 767 377 773 411
rect 807 377 813 411
rect 767 339 813 377
rect 767 305 773 339
rect 807 305 813 339
rect 767 267 813 305
rect 767 233 773 267
rect 807 233 813 267
rect 767 195 813 233
rect 767 161 773 195
rect 807 161 813 195
rect 767 118 813 161
rect 925 1275 971 1318
rect 925 1241 931 1275
rect 965 1241 971 1275
rect 925 1203 971 1241
rect 925 1169 931 1203
rect 965 1169 971 1203
rect 925 1131 971 1169
rect 925 1097 931 1131
rect 965 1097 971 1131
rect 925 1059 971 1097
rect 925 1025 931 1059
rect 965 1025 971 1059
rect 925 987 971 1025
rect 925 953 931 987
rect 965 953 971 987
rect 925 915 971 953
rect 925 881 931 915
rect 965 881 971 915
rect 925 843 971 881
rect 925 809 931 843
rect 965 809 971 843
rect 925 771 971 809
rect 925 737 931 771
rect 965 737 971 771
rect 925 699 971 737
rect 925 665 931 699
rect 965 665 971 699
rect 925 627 971 665
rect 925 593 931 627
rect 965 593 971 627
rect 925 555 971 593
rect 925 521 931 555
rect 965 521 971 555
rect 925 483 971 521
rect 925 449 931 483
rect 965 449 971 483
rect 925 411 971 449
rect 925 377 931 411
rect 965 377 971 411
rect 925 339 971 377
rect 925 305 931 339
rect 965 305 971 339
rect 925 267 971 305
rect 925 233 931 267
rect 965 233 971 267
rect 925 195 971 233
rect 925 161 931 195
rect 965 161 971 195
rect 925 118 971 161
rect 1083 1275 1129 1318
rect 1083 1241 1089 1275
rect 1123 1241 1129 1275
rect 1083 1203 1129 1241
rect 1083 1169 1089 1203
rect 1123 1169 1129 1203
rect 1083 1131 1129 1169
rect 1083 1097 1089 1131
rect 1123 1097 1129 1131
rect 1083 1059 1129 1097
rect 1083 1025 1089 1059
rect 1123 1025 1129 1059
rect 1083 987 1129 1025
rect 1083 953 1089 987
rect 1123 953 1129 987
rect 1083 915 1129 953
rect 1083 881 1089 915
rect 1123 881 1129 915
rect 1083 843 1129 881
rect 1083 809 1089 843
rect 1123 809 1129 843
rect 1083 771 1129 809
rect 1083 737 1089 771
rect 1123 737 1129 771
rect 1083 699 1129 737
rect 1083 665 1089 699
rect 1123 665 1129 699
rect 1083 627 1129 665
rect 1083 593 1089 627
rect 1123 593 1129 627
rect 1083 555 1129 593
rect 1083 521 1089 555
rect 1123 521 1129 555
rect 1083 483 1129 521
rect 1083 449 1089 483
rect 1123 449 1129 483
rect 1083 411 1129 449
rect 1083 377 1089 411
rect 1123 377 1129 411
rect 1083 339 1129 377
rect 1083 305 1089 339
rect 1123 305 1129 339
rect 1083 267 1129 305
rect 1083 233 1089 267
rect 1123 233 1129 267
rect 1083 195 1129 233
rect 1083 161 1089 195
rect 1123 161 1129 195
rect 1083 118 1129 161
rect -1073 71 -981 77
rect -1073 37 -1044 71
rect -1010 37 -981 71
rect -1073 31 -981 37
rect -915 71 -823 77
rect -915 37 -886 71
rect -852 37 -823 71
rect -915 31 -823 37
rect -757 71 -665 77
rect -757 37 -728 71
rect -694 37 -665 71
rect -757 31 -665 37
rect -599 71 -507 77
rect -599 37 -570 71
rect -536 37 -507 71
rect -599 31 -507 37
rect -441 71 -349 77
rect -441 37 -412 71
rect -378 37 -349 71
rect -441 31 -349 37
rect -283 71 -191 77
rect -283 37 -254 71
rect -220 37 -191 71
rect -283 31 -191 37
rect -125 71 -33 77
rect -125 37 -96 71
rect -62 37 -33 71
rect -125 31 -33 37
rect 33 71 125 77
rect 33 37 62 71
rect 96 37 125 71
rect 33 31 125 37
rect 191 71 283 77
rect 191 37 220 71
rect 254 37 283 71
rect 191 31 283 37
rect 349 71 441 77
rect 349 37 378 71
rect 412 37 441 71
rect 349 31 441 37
rect 507 71 599 77
rect 507 37 536 71
rect 570 37 599 71
rect 507 31 599 37
rect 665 71 757 77
rect 665 37 694 71
rect 728 37 757 71
rect 665 31 757 37
rect 823 71 915 77
rect 823 37 852 71
rect 886 37 915 71
rect 823 31 915 37
rect 981 71 1073 77
rect 981 37 1010 71
rect 1044 37 1073 71
rect 981 31 1073 37
rect -1129 -90 -1083 -47
rect -1129 -124 -1123 -90
rect -1089 -124 -1083 -90
rect -1129 -162 -1083 -124
rect -1129 -196 -1123 -162
rect -1089 -196 -1083 -162
rect -1129 -234 -1083 -196
rect -1129 -268 -1123 -234
rect -1089 -268 -1083 -234
rect -1129 -306 -1083 -268
rect -1129 -340 -1123 -306
rect -1089 -340 -1083 -306
rect -1129 -378 -1083 -340
rect -1129 -412 -1123 -378
rect -1089 -412 -1083 -378
rect -1129 -450 -1083 -412
rect -1129 -484 -1123 -450
rect -1089 -484 -1083 -450
rect -1129 -522 -1083 -484
rect -1129 -556 -1123 -522
rect -1089 -556 -1083 -522
rect -1129 -594 -1083 -556
rect -1129 -628 -1123 -594
rect -1089 -628 -1083 -594
rect -1129 -666 -1083 -628
rect -1129 -700 -1123 -666
rect -1089 -700 -1083 -666
rect -1129 -738 -1083 -700
rect -1129 -772 -1123 -738
rect -1089 -772 -1083 -738
rect -1129 -810 -1083 -772
rect -1129 -844 -1123 -810
rect -1089 -844 -1083 -810
rect -1129 -882 -1083 -844
rect -1129 -916 -1123 -882
rect -1089 -916 -1083 -882
rect -1129 -954 -1083 -916
rect -1129 -988 -1123 -954
rect -1089 -988 -1083 -954
rect -1129 -1026 -1083 -988
rect -1129 -1060 -1123 -1026
rect -1089 -1060 -1083 -1026
rect -1129 -1098 -1083 -1060
rect -1129 -1132 -1123 -1098
rect -1089 -1132 -1083 -1098
rect -1129 -1170 -1083 -1132
rect -1129 -1204 -1123 -1170
rect -1089 -1204 -1083 -1170
rect -1129 -1247 -1083 -1204
rect -971 -90 -925 -47
rect -971 -124 -965 -90
rect -931 -124 -925 -90
rect -971 -162 -925 -124
rect -971 -196 -965 -162
rect -931 -196 -925 -162
rect -971 -234 -925 -196
rect -971 -268 -965 -234
rect -931 -268 -925 -234
rect -971 -306 -925 -268
rect -971 -340 -965 -306
rect -931 -340 -925 -306
rect -971 -378 -925 -340
rect -971 -412 -965 -378
rect -931 -412 -925 -378
rect -971 -450 -925 -412
rect -971 -484 -965 -450
rect -931 -484 -925 -450
rect -971 -522 -925 -484
rect -971 -556 -965 -522
rect -931 -556 -925 -522
rect -971 -594 -925 -556
rect -971 -628 -965 -594
rect -931 -628 -925 -594
rect -971 -666 -925 -628
rect -971 -700 -965 -666
rect -931 -700 -925 -666
rect -971 -738 -925 -700
rect -971 -772 -965 -738
rect -931 -772 -925 -738
rect -971 -810 -925 -772
rect -971 -844 -965 -810
rect -931 -844 -925 -810
rect -971 -882 -925 -844
rect -971 -916 -965 -882
rect -931 -916 -925 -882
rect -971 -954 -925 -916
rect -971 -988 -965 -954
rect -931 -988 -925 -954
rect -971 -1026 -925 -988
rect -971 -1060 -965 -1026
rect -931 -1060 -925 -1026
rect -971 -1098 -925 -1060
rect -971 -1132 -965 -1098
rect -931 -1132 -925 -1098
rect -971 -1170 -925 -1132
rect -971 -1204 -965 -1170
rect -931 -1204 -925 -1170
rect -971 -1247 -925 -1204
rect -813 -90 -767 -47
rect -813 -124 -807 -90
rect -773 -124 -767 -90
rect -813 -162 -767 -124
rect -813 -196 -807 -162
rect -773 -196 -767 -162
rect -813 -234 -767 -196
rect -813 -268 -807 -234
rect -773 -268 -767 -234
rect -813 -306 -767 -268
rect -813 -340 -807 -306
rect -773 -340 -767 -306
rect -813 -378 -767 -340
rect -813 -412 -807 -378
rect -773 -412 -767 -378
rect -813 -450 -767 -412
rect -813 -484 -807 -450
rect -773 -484 -767 -450
rect -813 -522 -767 -484
rect -813 -556 -807 -522
rect -773 -556 -767 -522
rect -813 -594 -767 -556
rect -813 -628 -807 -594
rect -773 -628 -767 -594
rect -813 -666 -767 -628
rect -813 -700 -807 -666
rect -773 -700 -767 -666
rect -813 -738 -767 -700
rect -813 -772 -807 -738
rect -773 -772 -767 -738
rect -813 -810 -767 -772
rect -813 -844 -807 -810
rect -773 -844 -767 -810
rect -813 -882 -767 -844
rect -813 -916 -807 -882
rect -773 -916 -767 -882
rect -813 -954 -767 -916
rect -813 -988 -807 -954
rect -773 -988 -767 -954
rect -813 -1026 -767 -988
rect -813 -1060 -807 -1026
rect -773 -1060 -767 -1026
rect -813 -1098 -767 -1060
rect -813 -1132 -807 -1098
rect -773 -1132 -767 -1098
rect -813 -1170 -767 -1132
rect -813 -1204 -807 -1170
rect -773 -1204 -767 -1170
rect -813 -1247 -767 -1204
rect -655 -90 -609 -47
rect -655 -124 -649 -90
rect -615 -124 -609 -90
rect -655 -162 -609 -124
rect -655 -196 -649 -162
rect -615 -196 -609 -162
rect -655 -234 -609 -196
rect -655 -268 -649 -234
rect -615 -268 -609 -234
rect -655 -306 -609 -268
rect -655 -340 -649 -306
rect -615 -340 -609 -306
rect -655 -378 -609 -340
rect -655 -412 -649 -378
rect -615 -412 -609 -378
rect -655 -450 -609 -412
rect -655 -484 -649 -450
rect -615 -484 -609 -450
rect -655 -522 -609 -484
rect -655 -556 -649 -522
rect -615 -556 -609 -522
rect -655 -594 -609 -556
rect -655 -628 -649 -594
rect -615 -628 -609 -594
rect -655 -666 -609 -628
rect -655 -700 -649 -666
rect -615 -700 -609 -666
rect -655 -738 -609 -700
rect -655 -772 -649 -738
rect -615 -772 -609 -738
rect -655 -810 -609 -772
rect -655 -844 -649 -810
rect -615 -844 -609 -810
rect -655 -882 -609 -844
rect -655 -916 -649 -882
rect -615 -916 -609 -882
rect -655 -954 -609 -916
rect -655 -988 -649 -954
rect -615 -988 -609 -954
rect -655 -1026 -609 -988
rect -655 -1060 -649 -1026
rect -615 -1060 -609 -1026
rect -655 -1098 -609 -1060
rect -655 -1132 -649 -1098
rect -615 -1132 -609 -1098
rect -655 -1170 -609 -1132
rect -655 -1204 -649 -1170
rect -615 -1204 -609 -1170
rect -655 -1247 -609 -1204
rect -497 -90 -451 -47
rect -497 -124 -491 -90
rect -457 -124 -451 -90
rect -497 -162 -451 -124
rect -497 -196 -491 -162
rect -457 -196 -451 -162
rect -497 -234 -451 -196
rect -497 -268 -491 -234
rect -457 -268 -451 -234
rect -497 -306 -451 -268
rect -497 -340 -491 -306
rect -457 -340 -451 -306
rect -497 -378 -451 -340
rect -497 -412 -491 -378
rect -457 -412 -451 -378
rect -497 -450 -451 -412
rect -497 -484 -491 -450
rect -457 -484 -451 -450
rect -497 -522 -451 -484
rect -497 -556 -491 -522
rect -457 -556 -451 -522
rect -497 -594 -451 -556
rect -497 -628 -491 -594
rect -457 -628 -451 -594
rect -497 -666 -451 -628
rect -497 -700 -491 -666
rect -457 -700 -451 -666
rect -497 -738 -451 -700
rect -497 -772 -491 -738
rect -457 -772 -451 -738
rect -497 -810 -451 -772
rect -497 -844 -491 -810
rect -457 -844 -451 -810
rect -497 -882 -451 -844
rect -497 -916 -491 -882
rect -457 -916 -451 -882
rect -497 -954 -451 -916
rect -497 -988 -491 -954
rect -457 -988 -451 -954
rect -497 -1026 -451 -988
rect -497 -1060 -491 -1026
rect -457 -1060 -451 -1026
rect -497 -1098 -451 -1060
rect -497 -1132 -491 -1098
rect -457 -1132 -451 -1098
rect -497 -1170 -451 -1132
rect -497 -1204 -491 -1170
rect -457 -1204 -451 -1170
rect -497 -1247 -451 -1204
rect -339 -90 -293 -47
rect -339 -124 -333 -90
rect -299 -124 -293 -90
rect -339 -162 -293 -124
rect -339 -196 -333 -162
rect -299 -196 -293 -162
rect -339 -234 -293 -196
rect -339 -268 -333 -234
rect -299 -268 -293 -234
rect -339 -306 -293 -268
rect -339 -340 -333 -306
rect -299 -340 -293 -306
rect -339 -378 -293 -340
rect -339 -412 -333 -378
rect -299 -412 -293 -378
rect -339 -450 -293 -412
rect -339 -484 -333 -450
rect -299 -484 -293 -450
rect -339 -522 -293 -484
rect -339 -556 -333 -522
rect -299 -556 -293 -522
rect -339 -594 -293 -556
rect -339 -628 -333 -594
rect -299 -628 -293 -594
rect -339 -666 -293 -628
rect -339 -700 -333 -666
rect -299 -700 -293 -666
rect -339 -738 -293 -700
rect -339 -772 -333 -738
rect -299 -772 -293 -738
rect -339 -810 -293 -772
rect -339 -844 -333 -810
rect -299 -844 -293 -810
rect -339 -882 -293 -844
rect -339 -916 -333 -882
rect -299 -916 -293 -882
rect -339 -954 -293 -916
rect -339 -988 -333 -954
rect -299 -988 -293 -954
rect -339 -1026 -293 -988
rect -339 -1060 -333 -1026
rect -299 -1060 -293 -1026
rect -339 -1098 -293 -1060
rect -339 -1132 -333 -1098
rect -299 -1132 -293 -1098
rect -339 -1170 -293 -1132
rect -339 -1204 -333 -1170
rect -299 -1204 -293 -1170
rect -339 -1247 -293 -1204
rect -181 -90 -135 -47
rect -181 -124 -175 -90
rect -141 -124 -135 -90
rect -181 -162 -135 -124
rect -181 -196 -175 -162
rect -141 -196 -135 -162
rect -181 -234 -135 -196
rect -181 -268 -175 -234
rect -141 -268 -135 -234
rect -181 -306 -135 -268
rect -181 -340 -175 -306
rect -141 -340 -135 -306
rect -181 -378 -135 -340
rect -181 -412 -175 -378
rect -141 -412 -135 -378
rect -181 -450 -135 -412
rect -181 -484 -175 -450
rect -141 -484 -135 -450
rect -181 -522 -135 -484
rect -181 -556 -175 -522
rect -141 -556 -135 -522
rect -181 -594 -135 -556
rect -181 -628 -175 -594
rect -141 -628 -135 -594
rect -181 -666 -135 -628
rect -181 -700 -175 -666
rect -141 -700 -135 -666
rect -181 -738 -135 -700
rect -181 -772 -175 -738
rect -141 -772 -135 -738
rect -181 -810 -135 -772
rect -181 -844 -175 -810
rect -141 -844 -135 -810
rect -181 -882 -135 -844
rect -181 -916 -175 -882
rect -141 -916 -135 -882
rect -181 -954 -135 -916
rect -181 -988 -175 -954
rect -141 -988 -135 -954
rect -181 -1026 -135 -988
rect -181 -1060 -175 -1026
rect -141 -1060 -135 -1026
rect -181 -1098 -135 -1060
rect -181 -1132 -175 -1098
rect -141 -1132 -135 -1098
rect -181 -1170 -135 -1132
rect -181 -1204 -175 -1170
rect -141 -1204 -135 -1170
rect -181 -1247 -135 -1204
rect -23 -90 23 -47
rect -23 -124 -17 -90
rect 17 -124 23 -90
rect -23 -162 23 -124
rect -23 -196 -17 -162
rect 17 -196 23 -162
rect -23 -234 23 -196
rect -23 -268 -17 -234
rect 17 -268 23 -234
rect -23 -306 23 -268
rect -23 -340 -17 -306
rect 17 -340 23 -306
rect -23 -378 23 -340
rect -23 -412 -17 -378
rect 17 -412 23 -378
rect -23 -450 23 -412
rect -23 -484 -17 -450
rect 17 -484 23 -450
rect -23 -522 23 -484
rect -23 -556 -17 -522
rect 17 -556 23 -522
rect -23 -594 23 -556
rect -23 -628 -17 -594
rect 17 -628 23 -594
rect -23 -666 23 -628
rect -23 -700 -17 -666
rect 17 -700 23 -666
rect -23 -738 23 -700
rect -23 -772 -17 -738
rect 17 -772 23 -738
rect -23 -810 23 -772
rect -23 -844 -17 -810
rect 17 -844 23 -810
rect -23 -882 23 -844
rect -23 -916 -17 -882
rect 17 -916 23 -882
rect -23 -954 23 -916
rect -23 -988 -17 -954
rect 17 -988 23 -954
rect -23 -1026 23 -988
rect -23 -1060 -17 -1026
rect 17 -1060 23 -1026
rect -23 -1098 23 -1060
rect -23 -1132 -17 -1098
rect 17 -1132 23 -1098
rect -23 -1170 23 -1132
rect -23 -1204 -17 -1170
rect 17 -1204 23 -1170
rect -23 -1247 23 -1204
rect 135 -90 181 -47
rect 135 -124 141 -90
rect 175 -124 181 -90
rect 135 -162 181 -124
rect 135 -196 141 -162
rect 175 -196 181 -162
rect 135 -234 181 -196
rect 135 -268 141 -234
rect 175 -268 181 -234
rect 135 -306 181 -268
rect 135 -340 141 -306
rect 175 -340 181 -306
rect 135 -378 181 -340
rect 135 -412 141 -378
rect 175 -412 181 -378
rect 135 -450 181 -412
rect 135 -484 141 -450
rect 175 -484 181 -450
rect 135 -522 181 -484
rect 135 -556 141 -522
rect 175 -556 181 -522
rect 135 -594 181 -556
rect 135 -628 141 -594
rect 175 -628 181 -594
rect 135 -666 181 -628
rect 135 -700 141 -666
rect 175 -700 181 -666
rect 135 -738 181 -700
rect 135 -772 141 -738
rect 175 -772 181 -738
rect 135 -810 181 -772
rect 135 -844 141 -810
rect 175 -844 181 -810
rect 135 -882 181 -844
rect 135 -916 141 -882
rect 175 -916 181 -882
rect 135 -954 181 -916
rect 135 -988 141 -954
rect 175 -988 181 -954
rect 135 -1026 181 -988
rect 135 -1060 141 -1026
rect 175 -1060 181 -1026
rect 135 -1098 181 -1060
rect 135 -1132 141 -1098
rect 175 -1132 181 -1098
rect 135 -1170 181 -1132
rect 135 -1204 141 -1170
rect 175 -1204 181 -1170
rect 135 -1247 181 -1204
rect 293 -90 339 -47
rect 293 -124 299 -90
rect 333 -124 339 -90
rect 293 -162 339 -124
rect 293 -196 299 -162
rect 333 -196 339 -162
rect 293 -234 339 -196
rect 293 -268 299 -234
rect 333 -268 339 -234
rect 293 -306 339 -268
rect 293 -340 299 -306
rect 333 -340 339 -306
rect 293 -378 339 -340
rect 293 -412 299 -378
rect 333 -412 339 -378
rect 293 -450 339 -412
rect 293 -484 299 -450
rect 333 -484 339 -450
rect 293 -522 339 -484
rect 293 -556 299 -522
rect 333 -556 339 -522
rect 293 -594 339 -556
rect 293 -628 299 -594
rect 333 -628 339 -594
rect 293 -666 339 -628
rect 293 -700 299 -666
rect 333 -700 339 -666
rect 293 -738 339 -700
rect 293 -772 299 -738
rect 333 -772 339 -738
rect 293 -810 339 -772
rect 293 -844 299 -810
rect 333 -844 339 -810
rect 293 -882 339 -844
rect 293 -916 299 -882
rect 333 -916 339 -882
rect 293 -954 339 -916
rect 293 -988 299 -954
rect 333 -988 339 -954
rect 293 -1026 339 -988
rect 293 -1060 299 -1026
rect 333 -1060 339 -1026
rect 293 -1098 339 -1060
rect 293 -1132 299 -1098
rect 333 -1132 339 -1098
rect 293 -1170 339 -1132
rect 293 -1204 299 -1170
rect 333 -1204 339 -1170
rect 293 -1247 339 -1204
rect 451 -90 497 -47
rect 451 -124 457 -90
rect 491 -124 497 -90
rect 451 -162 497 -124
rect 451 -196 457 -162
rect 491 -196 497 -162
rect 451 -234 497 -196
rect 451 -268 457 -234
rect 491 -268 497 -234
rect 451 -306 497 -268
rect 451 -340 457 -306
rect 491 -340 497 -306
rect 451 -378 497 -340
rect 451 -412 457 -378
rect 491 -412 497 -378
rect 451 -450 497 -412
rect 451 -484 457 -450
rect 491 -484 497 -450
rect 451 -522 497 -484
rect 451 -556 457 -522
rect 491 -556 497 -522
rect 451 -594 497 -556
rect 451 -628 457 -594
rect 491 -628 497 -594
rect 451 -666 497 -628
rect 451 -700 457 -666
rect 491 -700 497 -666
rect 451 -738 497 -700
rect 451 -772 457 -738
rect 491 -772 497 -738
rect 451 -810 497 -772
rect 451 -844 457 -810
rect 491 -844 497 -810
rect 451 -882 497 -844
rect 451 -916 457 -882
rect 491 -916 497 -882
rect 451 -954 497 -916
rect 451 -988 457 -954
rect 491 -988 497 -954
rect 451 -1026 497 -988
rect 451 -1060 457 -1026
rect 491 -1060 497 -1026
rect 451 -1098 497 -1060
rect 451 -1132 457 -1098
rect 491 -1132 497 -1098
rect 451 -1170 497 -1132
rect 451 -1204 457 -1170
rect 491 -1204 497 -1170
rect 451 -1247 497 -1204
rect 609 -90 655 -47
rect 609 -124 615 -90
rect 649 -124 655 -90
rect 609 -162 655 -124
rect 609 -196 615 -162
rect 649 -196 655 -162
rect 609 -234 655 -196
rect 609 -268 615 -234
rect 649 -268 655 -234
rect 609 -306 655 -268
rect 609 -340 615 -306
rect 649 -340 655 -306
rect 609 -378 655 -340
rect 609 -412 615 -378
rect 649 -412 655 -378
rect 609 -450 655 -412
rect 609 -484 615 -450
rect 649 -484 655 -450
rect 609 -522 655 -484
rect 609 -556 615 -522
rect 649 -556 655 -522
rect 609 -594 655 -556
rect 609 -628 615 -594
rect 649 -628 655 -594
rect 609 -666 655 -628
rect 609 -700 615 -666
rect 649 -700 655 -666
rect 609 -738 655 -700
rect 609 -772 615 -738
rect 649 -772 655 -738
rect 609 -810 655 -772
rect 609 -844 615 -810
rect 649 -844 655 -810
rect 609 -882 655 -844
rect 609 -916 615 -882
rect 649 -916 655 -882
rect 609 -954 655 -916
rect 609 -988 615 -954
rect 649 -988 655 -954
rect 609 -1026 655 -988
rect 609 -1060 615 -1026
rect 649 -1060 655 -1026
rect 609 -1098 655 -1060
rect 609 -1132 615 -1098
rect 649 -1132 655 -1098
rect 609 -1170 655 -1132
rect 609 -1204 615 -1170
rect 649 -1204 655 -1170
rect 609 -1247 655 -1204
rect 767 -90 813 -47
rect 767 -124 773 -90
rect 807 -124 813 -90
rect 767 -162 813 -124
rect 767 -196 773 -162
rect 807 -196 813 -162
rect 767 -234 813 -196
rect 767 -268 773 -234
rect 807 -268 813 -234
rect 767 -306 813 -268
rect 767 -340 773 -306
rect 807 -340 813 -306
rect 767 -378 813 -340
rect 767 -412 773 -378
rect 807 -412 813 -378
rect 767 -450 813 -412
rect 767 -484 773 -450
rect 807 -484 813 -450
rect 767 -522 813 -484
rect 767 -556 773 -522
rect 807 -556 813 -522
rect 767 -594 813 -556
rect 767 -628 773 -594
rect 807 -628 813 -594
rect 767 -666 813 -628
rect 767 -700 773 -666
rect 807 -700 813 -666
rect 767 -738 813 -700
rect 767 -772 773 -738
rect 807 -772 813 -738
rect 767 -810 813 -772
rect 767 -844 773 -810
rect 807 -844 813 -810
rect 767 -882 813 -844
rect 767 -916 773 -882
rect 807 -916 813 -882
rect 767 -954 813 -916
rect 767 -988 773 -954
rect 807 -988 813 -954
rect 767 -1026 813 -988
rect 767 -1060 773 -1026
rect 807 -1060 813 -1026
rect 767 -1098 813 -1060
rect 767 -1132 773 -1098
rect 807 -1132 813 -1098
rect 767 -1170 813 -1132
rect 767 -1204 773 -1170
rect 807 -1204 813 -1170
rect 767 -1247 813 -1204
rect 925 -90 971 -47
rect 925 -124 931 -90
rect 965 -124 971 -90
rect 925 -162 971 -124
rect 925 -196 931 -162
rect 965 -196 971 -162
rect 925 -234 971 -196
rect 925 -268 931 -234
rect 965 -268 971 -234
rect 925 -306 971 -268
rect 925 -340 931 -306
rect 965 -340 971 -306
rect 925 -378 971 -340
rect 925 -412 931 -378
rect 965 -412 971 -378
rect 925 -450 971 -412
rect 925 -484 931 -450
rect 965 -484 971 -450
rect 925 -522 971 -484
rect 925 -556 931 -522
rect 965 -556 971 -522
rect 925 -594 971 -556
rect 925 -628 931 -594
rect 965 -628 971 -594
rect 925 -666 971 -628
rect 925 -700 931 -666
rect 965 -700 971 -666
rect 925 -738 971 -700
rect 925 -772 931 -738
rect 965 -772 971 -738
rect 925 -810 971 -772
rect 925 -844 931 -810
rect 965 -844 971 -810
rect 925 -882 971 -844
rect 925 -916 931 -882
rect 965 -916 971 -882
rect 925 -954 971 -916
rect 925 -988 931 -954
rect 965 -988 971 -954
rect 925 -1026 971 -988
rect 925 -1060 931 -1026
rect 965 -1060 971 -1026
rect 925 -1098 971 -1060
rect 925 -1132 931 -1098
rect 965 -1132 971 -1098
rect 925 -1170 971 -1132
rect 925 -1204 931 -1170
rect 965 -1204 971 -1170
rect 925 -1247 971 -1204
rect 1083 -90 1129 -47
rect 1083 -124 1089 -90
rect 1123 -124 1129 -90
rect 1083 -162 1129 -124
rect 1083 -196 1089 -162
rect 1123 -196 1129 -162
rect 1083 -234 1129 -196
rect 1083 -268 1089 -234
rect 1123 -268 1129 -234
rect 1083 -306 1129 -268
rect 1083 -340 1089 -306
rect 1123 -340 1129 -306
rect 1083 -378 1129 -340
rect 1083 -412 1089 -378
rect 1123 -412 1129 -378
rect 1083 -450 1129 -412
rect 1083 -484 1089 -450
rect 1123 -484 1129 -450
rect 1083 -522 1129 -484
rect 1083 -556 1089 -522
rect 1123 -556 1129 -522
rect 1083 -594 1129 -556
rect 1083 -628 1089 -594
rect 1123 -628 1129 -594
rect 1083 -666 1129 -628
rect 1083 -700 1089 -666
rect 1123 -700 1129 -666
rect 1083 -738 1129 -700
rect 1083 -772 1089 -738
rect 1123 -772 1129 -738
rect 1083 -810 1129 -772
rect 1083 -844 1089 -810
rect 1123 -844 1129 -810
rect 1083 -882 1129 -844
rect 1083 -916 1089 -882
rect 1123 -916 1129 -882
rect 1083 -954 1129 -916
rect 1083 -988 1089 -954
rect 1123 -988 1129 -954
rect 1083 -1026 1129 -988
rect 1083 -1060 1089 -1026
rect 1123 -1060 1129 -1026
rect 1083 -1098 1129 -1060
rect 1083 -1132 1089 -1098
rect 1123 -1132 1129 -1098
rect 1083 -1170 1129 -1132
rect 1083 -1204 1089 -1170
rect 1123 -1204 1129 -1170
rect 1083 -1247 1129 -1204
rect -1073 -1294 -981 -1288
rect -1073 -1328 -1044 -1294
rect -1010 -1328 -981 -1294
rect -1073 -1334 -981 -1328
rect -915 -1294 -823 -1288
rect -915 -1328 -886 -1294
rect -852 -1328 -823 -1294
rect -915 -1334 -823 -1328
rect -757 -1294 -665 -1288
rect -757 -1328 -728 -1294
rect -694 -1328 -665 -1294
rect -757 -1334 -665 -1328
rect -599 -1294 -507 -1288
rect -599 -1328 -570 -1294
rect -536 -1328 -507 -1294
rect -599 -1334 -507 -1328
rect -441 -1294 -349 -1288
rect -441 -1328 -412 -1294
rect -378 -1328 -349 -1294
rect -441 -1334 -349 -1328
rect -283 -1294 -191 -1288
rect -283 -1328 -254 -1294
rect -220 -1328 -191 -1294
rect -283 -1334 -191 -1328
rect -125 -1294 -33 -1288
rect -125 -1328 -96 -1294
rect -62 -1328 -33 -1294
rect -125 -1334 -33 -1328
rect 33 -1294 125 -1288
rect 33 -1328 62 -1294
rect 96 -1328 125 -1294
rect 33 -1334 125 -1328
rect 191 -1294 283 -1288
rect 191 -1328 220 -1294
rect 254 -1328 283 -1294
rect 191 -1334 283 -1328
rect 349 -1294 441 -1288
rect 349 -1328 378 -1294
rect 412 -1328 441 -1294
rect 349 -1334 441 -1328
rect 507 -1294 599 -1288
rect 507 -1328 536 -1294
rect 570 -1328 599 -1294
rect 507 -1334 599 -1328
rect 665 -1294 757 -1288
rect 665 -1328 694 -1294
rect 728 -1328 757 -1294
rect 665 -1334 757 -1328
rect 823 -1294 915 -1288
rect 823 -1328 852 -1294
rect 886 -1328 915 -1294
rect 823 -1334 915 -1328
rect 981 -1294 1073 -1288
rect 981 -1328 1010 -1294
rect 1044 -1328 1073 -1294
rect 981 -1334 1073 -1328
rect -1129 -1455 -1083 -1412
rect -1129 -1489 -1123 -1455
rect -1089 -1489 -1083 -1455
rect -1129 -1527 -1083 -1489
rect -1129 -1561 -1123 -1527
rect -1089 -1561 -1083 -1527
rect -1129 -1599 -1083 -1561
rect -1129 -1633 -1123 -1599
rect -1089 -1633 -1083 -1599
rect -1129 -1671 -1083 -1633
rect -1129 -1705 -1123 -1671
rect -1089 -1705 -1083 -1671
rect -1129 -1743 -1083 -1705
rect -1129 -1777 -1123 -1743
rect -1089 -1777 -1083 -1743
rect -1129 -1815 -1083 -1777
rect -1129 -1849 -1123 -1815
rect -1089 -1849 -1083 -1815
rect -1129 -1887 -1083 -1849
rect -1129 -1921 -1123 -1887
rect -1089 -1921 -1083 -1887
rect -1129 -1959 -1083 -1921
rect -1129 -1993 -1123 -1959
rect -1089 -1993 -1083 -1959
rect -1129 -2031 -1083 -1993
rect -1129 -2065 -1123 -2031
rect -1089 -2065 -1083 -2031
rect -1129 -2103 -1083 -2065
rect -1129 -2137 -1123 -2103
rect -1089 -2137 -1083 -2103
rect -1129 -2175 -1083 -2137
rect -1129 -2209 -1123 -2175
rect -1089 -2209 -1083 -2175
rect -1129 -2247 -1083 -2209
rect -1129 -2281 -1123 -2247
rect -1089 -2281 -1083 -2247
rect -1129 -2319 -1083 -2281
rect -1129 -2353 -1123 -2319
rect -1089 -2353 -1083 -2319
rect -1129 -2391 -1083 -2353
rect -1129 -2425 -1123 -2391
rect -1089 -2425 -1083 -2391
rect -1129 -2463 -1083 -2425
rect -1129 -2497 -1123 -2463
rect -1089 -2497 -1083 -2463
rect -1129 -2535 -1083 -2497
rect -1129 -2569 -1123 -2535
rect -1089 -2569 -1083 -2535
rect -1129 -2612 -1083 -2569
rect -971 -1455 -925 -1412
rect -971 -1489 -965 -1455
rect -931 -1489 -925 -1455
rect -971 -1527 -925 -1489
rect -971 -1561 -965 -1527
rect -931 -1561 -925 -1527
rect -971 -1599 -925 -1561
rect -971 -1633 -965 -1599
rect -931 -1633 -925 -1599
rect -971 -1671 -925 -1633
rect -971 -1705 -965 -1671
rect -931 -1705 -925 -1671
rect -971 -1743 -925 -1705
rect -971 -1777 -965 -1743
rect -931 -1777 -925 -1743
rect -971 -1815 -925 -1777
rect -971 -1849 -965 -1815
rect -931 -1849 -925 -1815
rect -971 -1887 -925 -1849
rect -971 -1921 -965 -1887
rect -931 -1921 -925 -1887
rect -971 -1959 -925 -1921
rect -971 -1993 -965 -1959
rect -931 -1993 -925 -1959
rect -971 -2031 -925 -1993
rect -971 -2065 -965 -2031
rect -931 -2065 -925 -2031
rect -971 -2103 -925 -2065
rect -971 -2137 -965 -2103
rect -931 -2137 -925 -2103
rect -971 -2175 -925 -2137
rect -971 -2209 -965 -2175
rect -931 -2209 -925 -2175
rect -971 -2247 -925 -2209
rect -971 -2281 -965 -2247
rect -931 -2281 -925 -2247
rect -971 -2319 -925 -2281
rect -971 -2353 -965 -2319
rect -931 -2353 -925 -2319
rect -971 -2391 -925 -2353
rect -971 -2425 -965 -2391
rect -931 -2425 -925 -2391
rect -971 -2463 -925 -2425
rect -971 -2497 -965 -2463
rect -931 -2497 -925 -2463
rect -971 -2535 -925 -2497
rect -971 -2569 -965 -2535
rect -931 -2569 -925 -2535
rect -971 -2612 -925 -2569
rect -813 -1455 -767 -1412
rect -813 -1489 -807 -1455
rect -773 -1489 -767 -1455
rect -813 -1527 -767 -1489
rect -813 -1561 -807 -1527
rect -773 -1561 -767 -1527
rect -813 -1599 -767 -1561
rect -813 -1633 -807 -1599
rect -773 -1633 -767 -1599
rect -813 -1671 -767 -1633
rect -813 -1705 -807 -1671
rect -773 -1705 -767 -1671
rect -813 -1743 -767 -1705
rect -813 -1777 -807 -1743
rect -773 -1777 -767 -1743
rect -813 -1815 -767 -1777
rect -813 -1849 -807 -1815
rect -773 -1849 -767 -1815
rect -813 -1887 -767 -1849
rect -813 -1921 -807 -1887
rect -773 -1921 -767 -1887
rect -813 -1959 -767 -1921
rect -813 -1993 -807 -1959
rect -773 -1993 -767 -1959
rect -813 -2031 -767 -1993
rect -813 -2065 -807 -2031
rect -773 -2065 -767 -2031
rect -813 -2103 -767 -2065
rect -813 -2137 -807 -2103
rect -773 -2137 -767 -2103
rect -813 -2175 -767 -2137
rect -813 -2209 -807 -2175
rect -773 -2209 -767 -2175
rect -813 -2247 -767 -2209
rect -813 -2281 -807 -2247
rect -773 -2281 -767 -2247
rect -813 -2319 -767 -2281
rect -813 -2353 -807 -2319
rect -773 -2353 -767 -2319
rect -813 -2391 -767 -2353
rect -813 -2425 -807 -2391
rect -773 -2425 -767 -2391
rect -813 -2463 -767 -2425
rect -813 -2497 -807 -2463
rect -773 -2497 -767 -2463
rect -813 -2535 -767 -2497
rect -813 -2569 -807 -2535
rect -773 -2569 -767 -2535
rect -813 -2612 -767 -2569
rect -655 -1455 -609 -1412
rect -655 -1489 -649 -1455
rect -615 -1489 -609 -1455
rect -655 -1527 -609 -1489
rect -655 -1561 -649 -1527
rect -615 -1561 -609 -1527
rect -655 -1599 -609 -1561
rect -655 -1633 -649 -1599
rect -615 -1633 -609 -1599
rect -655 -1671 -609 -1633
rect -655 -1705 -649 -1671
rect -615 -1705 -609 -1671
rect -655 -1743 -609 -1705
rect -655 -1777 -649 -1743
rect -615 -1777 -609 -1743
rect -655 -1815 -609 -1777
rect -655 -1849 -649 -1815
rect -615 -1849 -609 -1815
rect -655 -1887 -609 -1849
rect -655 -1921 -649 -1887
rect -615 -1921 -609 -1887
rect -655 -1959 -609 -1921
rect -655 -1993 -649 -1959
rect -615 -1993 -609 -1959
rect -655 -2031 -609 -1993
rect -655 -2065 -649 -2031
rect -615 -2065 -609 -2031
rect -655 -2103 -609 -2065
rect -655 -2137 -649 -2103
rect -615 -2137 -609 -2103
rect -655 -2175 -609 -2137
rect -655 -2209 -649 -2175
rect -615 -2209 -609 -2175
rect -655 -2247 -609 -2209
rect -655 -2281 -649 -2247
rect -615 -2281 -609 -2247
rect -655 -2319 -609 -2281
rect -655 -2353 -649 -2319
rect -615 -2353 -609 -2319
rect -655 -2391 -609 -2353
rect -655 -2425 -649 -2391
rect -615 -2425 -609 -2391
rect -655 -2463 -609 -2425
rect -655 -2497 -649 -2463
rect -615 -2497 -609 -2463
rect -655 -2535 -609 -2497
rect -655 -2569 -649 -2535
rect -615 -2569 -609 -2535
rect -655 -2612 -609 -2569
rect -497 -1455 -451 -1412
rect -497 -1489 -491 -1455
rect -457 -1489 -451 -1455
rect -497 -1527 -451 -1489
rect -497 -1561 -491 -1527
rect -457 -1561 -451 -1527
rect -497 -1599 -451 -1561
rect -497 -1633 -491 -1599
rect -457 -1633 -451 -1599
rect -497 -1671 -451 -1633
rect -497 -1705 -491 -1671
rect -457 -1705 -451 -1671
rect -497 -1743 -451 -1705
rect -497 -1777 -491 -1743
rect -457 -1777 -451 -1743
rect -497 -1815 -451 -1777
rect -497 -1849 -491 -1815
rect -457 -1849 -451 -1815
rect -497 -1887 -451 -1849
rect -497 -1921 -491 -1887
rect -457 -1921 -451 -1887
rect -497 -1959 -451 -1921
rect -497 -1993 -491 -1959
rect -457 -1993 -451 -1959
rect -497 -2031 -451 -1993
rect -497 -2065 -491 -2031
rect -457 -2065 -451 -2031
rect -497 -2103 -451 -2065
rect -497 -2137 -491 -2103
rect -457 -2137 -451 -2103
rect -497 -2175 -451 -2137
rect -497 -2209 -491 -2175
rect -457 -2209 -451 -2175
rect -497 -2247 -451 -2209
rect -497 -2281 -491 -2247
rect -457 -2281 -451 -2247
rect -497 -2319 -451 -2281
rect -497 -2353 -491 -2319
rect -457 -2353 -451 -2319
rect -497 -2391 -451 -2353
rect -497 -2425 -491 -2391
rect -457 -2425 -451 -2391
rect -497 -2463 -451 -2425
rect -497 -2497 -491 -2463
rect -457 -2497 -451 -2463
rect -497 -2535 -451 -2497
rect -497 -2569 -491 -2535
rect -457 -2569 -451 -2535
rect -497 -2612 -451 -2569
rect -339 -1455 -293 -1412
rect -339 -1489 -333 -1455
rect -299 -1489 -293 -1455
rect -339 -1527 -293 -1489
rect -339 -1561 -333 -1527
rect -299 -1561 -293 -1527
rect -339 -1599 -293 -1561
rect -339 -1633 -333 -1599
rect -299 -1633 -293 -1599
rect -339 -1671 -293 -1633
rect -339 -1705 -333 -1671
rect -299 -1705 -293 -1671
rect -339 -1743 -293 -1705
rect -339 -1777 -333 -1743
rect -299 -1777 -293 -1743
rect -339 -1815 -293 -1777
rect -339 -1849 -333 -1815
rect -299 -1849 -293 -1815
rect -339 -1887 -293 -1849
rect -339 -1921 -333 -1887
rect -299 -1921 -293 -1887
rect -339 -1959 -293 -1921
rect -339 -1993 -333 -1959
rect -299 -1993 -293 -1959
rect -339 -2031 -293 -1993
rect -339 -2065 -333 -2031
rect -299 -2065 -293 -2031
rect -339 -2103 -293 -2065
rect -339 -2137 -333 -2103
rect -299 -2137 -293 -2103
rect -339 -2175 -293 -2137
rect -339 -2209 -333 -2175
rect -299 -2209 -293 -2175
rect -339 -2247 -293 -2209
rect -339 -2281 -333 -2247
rect -299 -2281 -293 -2247
rect -339 -2319 -293 -2281
rect -339 -2353 -333 -2319
rect -299 -2353 -293 -2319
rect -339 -2391 -293 -2353
rect -339 -2425 -333 -2391
rect -299 -2425 -293 -2391
rect -339 -2463 -293 -2425
rect -339 -2497 -333 -2463
rect -299 -2497 -293 -2463
rect -339 -2535 -293 -2497
rect -339 -2569 -333 -2535
rect -299 -2569 -293 -2535
rect -339 -2612 -293 -2569
rect -181 -1455 -135 -1412
rect -181 -1489 -175 -1455
rect -141 -1489 -135 -1455
rect -181 -1527 -135 -1489
rect -181 -1561 -175 -1527
rect -141 -1561 -135 -1527
rect -181 -1599 -135 -1561
rect -181 -1633 -175 -1599
rect -141 -1633 -135 -1599
rect -181 -1671 -135 -1633
rect -181 -1705 -175 -1671
rect -141 -1705 -135 -1671
rect -181 -1743 -135 -1705
rect -181 -1777 -175 -1743
rect -141 -1777 -135 -1743
rect -181 -1815 -135 -1777
rect -181 -1849 -175 -1815
rect -141 -1849 -135 -1815
rect -181 -1887 -135 -1849
rect -181 -1921 -175 -1887
rect -141 -1921 -135 -1887
rect -181 -1959 -135 -1921
rect -181 -1993 -175 -1959
rect -141 -1993 -135 -1959
rect -181 -2031 -135 -1993
rect -181 -2065 -175 -2031
rect -141 -2065 -135 -2031
rect -181 -2103 -135 -2065
rect -181 -2137 -175 -2103
rect -141 -2137 -135 -2103
rect -181 -2175 -135 -2137
rect -181 -2209 -175 -2175
rect -141 -2209 -135 -2175
rect -181 -2247 -135 -2209
rect -181 -2281 -175 -2247
rect -141 -2281 -135 -2247
rect -181 -2319 -135 -2281
rect -181 -2353 -175 -2319
rect -141 -2353 -135 -2319
rect -181 -2391 -135 -2353
rect -181 -2425 -175 -2391
rect -141 -2425 -135 -2391
rect -181 -2463 -135 -2425
rect -181 -2497 -175 -2463
rect -141 -2497 -135 -2463
rect -181 -2535 -135 -2497
rect -181 -2569 -175 -2535
rect -141 -2569 -135 -2535
rect -181 -2612 -135 -2569
rect -23 -1455 23 -1412
rect -23 -1489 -17 -1455
rect 17 -1489 23 -1455
rect -23 -1527 23 -1489
rect -23 -1561 -17 -1527
rect 17 -1561 23 -1527
rect -23 -1599 23 -1561
rect -23 -1633 -17 -1599
rect 17 -1633 23 -1599
rect -23 -1671 23 -1633
rect -23 -1705 -17 -1671
rect 17 -1705 23 -1671
rect -23 -1743 23 -1705
rect -23 -1777 -17 -1743
rect 17 -1777 23 -1743
rect -23 -1815 23 -1777
rect -23 -1849 -17 -1815
rect 17 -1849 23 -1815
rect -23 -1887 23 -1849
rect -23 -1921 -17 -1887
rect 17 -1921 23 -1887
rect -23 -1959 23 -1921
rect -23 -1993 -17 -1959
rect 17 -1993 23 -1959
rect -23 -2031 23 -1993
rect -23 -2065 -17 -2031
rect 17 -2065 23 -2031
rect -23 -2103 23 -2065
rect -23 -2137 -17 -2103
rect 17 -2137 23 -2103
rect -23 -2175 23 -2137
rect -23 -2209 -17 -2175
rect 17 -2209 23 -2175
rect -23 -2247 23 -2209
rect -23 -2281 -17 -2247
rect 17 -2281 23 -2247
rect -23 -2319 23 -2281
rect -23 -2353 -17 -2319
rect 17 -2353 23 -2319
rect -23 -2391 23 -2353
rect -23 -2425 -17 -2391
rect 17 -2425 23 -2391
rect -23 -2463 23 -2425
rect -23 -2497 -17 -2463
rect 17 -2497 23 -2463
rect -23 -2535 23 -2497
rect -23 -2569 -17 -2535
rect 17 -2569 23 -2535
rect -23 -2612 23 -2569
rect 135 -1455 181 -1412
rect 135 -1489 141 -1455
rect 175 -1489 181 -1455
rect 135 -1527 181 -1489
rect 135 -1561 141 -1527
rect 175 -1561 181 -1527
rect 135 -1599 181 -1561
rect 135 -1633 141 -1599
rect 175 -1633 181 -1599
rect 135 -1671 181 -1633
rect 135 -1705 141 -1671
rect 175 -1705 181 -1671
rect 135 -1743 181 -1705
rect 135 -1777 141 -1743
rect 175 -1777 181 -1743
rect 135 -1815 181 -1777
rect 135 -1849 141 -1815
rect 175 -1849 181 -1815
rect 135 -1887 181 -1849
rect 135 -1921 141 -1887
rect 175 -1921 181 -1887
rect 135 -1959 181 -1921
rect 135 -1993 141 -1959
rect 175 -1993 181 -1959
rect 135 -2031 181 -1993
rect 135 -2065 141 -2031
rect 175 -2065 181 -2031
rect 135 -2103 181 -2065
rect 135 -2137 141 -2103
rect 175 -2137 181 -2103
rect 135 -2175 181 -2137
rect 135 -2209 141 -2175
rect 175 -2209 181 -2175
rect 135 -2247 181 -2209
rect 135 -2281 141 -2247
rect 175 -2281 181 -2247
rect 135 -2319 181 -2281
rect 135 -2353 141 -2319
rect 175 -2353 181 -2319
rect 135 -2391 181 -2353
rect 135 -2425 141 -2391
rect 175 -2425 181 -2391
rect 135 -2463 181 -2425
rect 135 -2497 141 -2463
rect 175 -2497 181 -2463
rect 135 -2535 181 -2497
rect 135 -2569 141 -2535
rect 175 -2569 181 -2535
rect 135 -2612 181 -2569
rect 293 -1455 339 -1412
rect 293 -1489 299 -1455
rect 333 -1489 339 -1455
rect 293 -1527 339 -1489
rect 293 -1561 299 -1527
rect 333 -1561 339 -1527
rect 293 -1599 339 -1561
rect 293 -1633 299 -1599
rect 333 -1633 339 -1599
rect 293 -1671 339 -1633
rect 293 -1705 299 -1671
rect 333 -1705 339 -1671
rect 293 -1743 339 -1705
rect 293 -1777 299 -1743
rect 333 -1777 339 -1743
rect 293 -1815 339 -1777
rect 293 -1849 299 -1815
rect 333 -1849 339 -1815
rect 293 -1887 339 -1849
rect 293 -1921 299 -1887
rect 333 -1921 339 -1887
rect 293 -1959 339 -1921
rect 293 -1993 299 -1959
rect 333 -1993 339 -1959
rect 293 -2031 339 -1993
rect 293 -2065 299 -2031
rect 333 -2065 339 -2031
rect 293 -2103 339 -2065
rect 293 -2137 299 -2103
rect 333 -2137 339 -2103
rect 293 -2175 339 -2137
rect 293 -2209 299 -2175
rect 333 -2209 339 -2175
rect 293 -2247 339 -2209
rect 293 -2281 299 -2247
rect 333 -2281 339 -2247
rect 293 -2319 339 -2281
rect 293 -2353 299 -2319
rect 333 -2353 339 -2319
rect 293 -2391 339 -2353
rect 293 -2425 299 -2391
rect 333 -2425 339 -2391
rect 293 -2463 339 -2425
rect 293 -2497 299 -2463
rect 333 -2497 339 -2463
rect 293 -2535 339 -2497
rect 293 -2569 299 -2535
rect 333 -2569 339 -2535
rect 293 -2612 339 -2569
rect 451 -1455 497 -1412
rect 451 -1489 457 -1455
rect 491 -1489 497 -1455
rect 451 -1527 497 -1489
rect 451 -1561 457 -1527
rect 491 -1561 497 -1527
rect 451 -1599 497 -1561
rect 451 -1633 457 -1599
rect 491 -1633 497 -1599
rect 451 -1671 497 -1633
rect 451 -1705 457 -1671
rect 491 -1705 497 -1671
rect 451 -1743 497 -1705
rect 451 -1777 457 -1743
rect 491 -1777 497 -1743
rect 451 -1815 497 -1777
rect 451 -1849 457 -1815
rect 491 -1849 497 -1815
rect 451 -1887 497 -1849
rect 451 -1921 457 -1887
rect 491 -1921 497 -1887
rect 451 -1959 497 -1921
rect 451 -1993 457 -1959
rect 491 -1993 497 -1959
rect 451 -2031 497 -1993
rect 451 -2065 457 -2031
rect 491 -2065 497 -2031
rect 451 -2103 497 -2065
rect 451 -2137 457 -2103
rect 491 -2137 497 -2103
rect 451 -2175 497 -2137
rect 451 -2209 457 -2175
rect 491 -2209 497 -2175
rect 451 -2247 497 -2209
rect 451 -2281 457 -2247
rect 491 -2281 497 -2247
rect 451 -2319 497 -2281
rect 451 -2353 457 -2319
rect 491 -2353 497 -2319
rect 451 -2391 497 -2353
rect 451 -2425 457 -2391
rect 491 -2425 497 -2391
rect 451 -2463 497 -2425
rect 451 -2497 457 -2463
rect 491 -2497 497 -2463
rect 451 -2535 497 -2497
rect 451 -2569 457 -2535
rect 491 -2569 497 -2535
rect 451 -2612 497 -2569
rect 609 -1455 655 -1412
rect 609 -1489 615 -1455
rect 649 -1489 655 -1455
rect 609 -1527 655 -1489
rect 609 -1561 615 -1527
rect 649 -1561 655 -1527
rect 609 -1599 655 -1561
rect 609 -1633 615 -1599
rect 649 -1633 655 -1599
rect 609 -1671 655 -1633
rect 609 -1705 615 -1671
rect 649 -1705 655 -1671
rect 609 -1743 655 -1705
rect 609 -1777 615 -1743
rect 649 -1777 655 -1743
rect 609 -1815 655 -1777
rect 609 -1849 615 -1815
rect 649 -1849 655 -1815
rect 609 -1887 655 -1849
rect 609 -1921 615 -1887
rect 649 -1921 655 -1887
rect 609 -1959 655 -1921
rect 609 -1993 615 -1959
rect 649 -1993 655 -1959
rect 609 -2031 655 -1993
rect 609 -2065 615 -2031
rect 649 -2065 655 -2031
rect 609 -2103 655 -2065
rect 609 -2137 615 -2103
rect 649 -2137 655 -2103
rect 609 -2175 655 -2137
rect 609 -2209 615 -2175
rect 649 -2209 655 -2175
rect 609 -2247 655 -2209
rect 609 -2281 615 -2247
rect 649 -2281 655 -2247
rect 609 -2319 655 -2281
rect 609 -2353 615 -2319
rect 649 -2353 655 -2319
rect 609 -2391 655 -2353
rect 609 -2425 615 -2391
rect 649 -2425 655 -2391
rect 609 -2463 655 -2425
rect 609 -2497 615 -2463
rect 649 -2497 655 -2463
rect 609 -2535 655 -2497
rect 609 -2569 615 -2535
rect 649 -2569 655 -2535
rect 609 -2612 655 -2569
rect 767 -1455 813 -1412
rect 767 -1489 773 -1455
rect 807 -1489 813 -1455
rect 767 -1527 813 -1489
rect 767 -1561 773 -1527
rect 807 -1561 813 -1527
rect 767 -1599 813 -1561
rect 767 -1633 773 -1599
rect 807 -1633 813 -1599
rect 767 -1671 813 -1633
rect 767 -1705 773 -1671
rect 807 -1705 813 -1671
rect 767 -1743 813 -1705
rect 767 -1777 773 -1743
rect 807 -1777 813 -1743
rect 767 -1815 813 -1777
rect 767 -1849 773 -1815
rect 807 -1849 813 -1815
rect 767 -1887 813 -1849
rect 767 -1921 773 -1887
rect 807 -1921 813 -1887
rect 767 -1959 813 -1921
rect 767 -1993 773 -1959
rect 807 -1993 813 -1959
rect 767 -2031 813 -1993
rect 767 -2065 773 -2031
rect 807 -2065 813 -2031
rect 767 -2103 813 -2065
rect 767 -2137 773 -2103
rect 807 -2137 813 -2103
rect 767 -2175 813 -2137
rect 767 -2209 773 -2175
rect 807 -2209 813 -2175
rect 767 -2247 813 -2209
rect 767 -2281 773 -2247
rect 807 -2281 813 -2247
rect 767 -2319 813 -2281
rect 767 -2353 773 -2319
rect 807 -2353 813 -2319
rect 767 -2391 813 -2353
rect 767 -2425 773 -2391
rect 807 -2425 813 -2391
rect 767 -2463 813 -2425
rect 767 -2497 773 -2463
rect 807 -2497 813 -2463
rect 767 -2535 813 -2497
rect 767 -2569 773 -2535
rect 807 -2569 813 -2535
rect 767 -2612 813 -2569
rect 925 -1455 971 -1412
rect 925 -1489 931 -1455
rect 965 -1489 971 -1455
rect 925 -1527 971 -1489
rect 925 -1561 931 -1527
rect 965 -1561 971 -1527
rect 925 -1599 971 -1561
rect 925 -1633 931 -1599
rect 965 -1633 971 -1599
rect 925 -1671 971 -1633
rect 925 -1705 931 -1671
rect 965 -1705 971 -1671
rect 925 -1743 971 -1705
rect 925 -1777 931 -1743
rect 965 -1777 971 -1743
rect 925 -1815 971 -1777
rect 925 -1849 931 -1815
rect 965 -1849 971 -1815
rect 925 -1887 971 -1849
rect 925 -1921 931 -1887
rect 965 -1921 971 -1887
rect 925 -1959 971 -1921
rect 925 -1993 931 -1959
rect 965 -1993 971 -1959
rect 925 -2031 971 -1993
rect 925 -2065 931 -2031
rect 965 -2065 971 -2031
rect 925 -2103 971 -2065
rect 925 -2137 931 -2103
rect 965 -2137 971 -2103
rect 925 -2175 971 -2137
rect 925 -2209 931 -2175
rect 965 -2209 971 -2175
rect 925 -2247 971 -2209
rect 925 -2281 931 -2247
rect 965 -2281 971 -2247
rect 925 -2319 971 -2281
rect 925 -2353 931 -2319
rect 965 -2353 971 -2319
rect 925 -2391 971 -2353
rect 925 -2425 931 -2391
rect 965 -2425 971 -2391
rect 925 -2463 971 -2425
rect 925 -2497 931 -2463
rect 965 -2497 971 -2463
rect 925 -2535 971 -2497
rect 925 -2569 931 -2535
rect 965 -2569 971 -2535
rect 925 -2612 971 -2569
rect 1083 -1455 1129 -1412
rect 1083 -1489 1089 -1455
rect 1123 -1489 1129 -1455
rect 1083 -1527 1129 -1489
rect 1083 -1561 1089 -1527
rect 1123 -1561 1129 -1527
rect 1083 -1599 1129 -1561
rect 1083 -1633 1089 -1599
rect 1123 -1633 1129 -1599
rect 1083 -1671 1129 -1633
rect 1083 -1705 1089 -1671
rect 1123 -1705 1129 -1671
rect 1083 -1743 1129 -1705
rect 1083 -1777 1089 -1743
rect 1123 -1777 1129 -1743
rect 1083 -1815 1129 -1777
rect 1083 -1849 1089 -1815
rect 1123 -1849 1129 -1815
rect 1083 -1887 1129 -1849
rect 1083 -1921 1089 -1887
rect 1123 -1921 1129 -1887
rect 1083 -1959 1129 -1921
rect 1083 -1993 1089 -1959
rect 1123 -1993 1129 -1959
rect 1083 -2031 1129 -1993
rect 1083 -2065 1089 -2031
rect 1123 -2065 1129 -2031
rect 1083 -2103 1129 -2065
rect 1083 -2137 1089 -2103
rect 1123 -2137 1129 -2103
rect 1083 -2175 1129 -2137
rect 1083 -2209 1089 -2175
rect 1123 -2209 1129 -2175
rect 1083 -2247 1129 -2209
rect 1083 -2281 1089 -2247
rect 1123 -2281 1129 -2247
rect 1083 -2319 1129 -2281
rect 1083 -2353 1089 -2319
rect 1123 -2353 1129 -2319
rect 1083 -2391 1129 -2353
rect 1083 -2425 1089 -2391
rect 1123 -2425 1129 -2391
rect 1083 -2463 1129 -2425
rect 1083 -2497 1089 -2463
rect 1123 -2497 1129 -2463
rect 1083 -2535 1129 -2497
rect 1083 -2569 1089 -2535
rect 1123 -2569 1129 -2535
rect 1083 -2612 1129 -2569
rect -1073 -2659 -981 -2653
rect -1073 -2693 -1044 -2659
rect -1010 -2693 -981 -2659
rect -1073 -2699 -981 -2693
rect -915 -2659 -823 -2653
rect -915 -2693 -886 -2659
rect -852 -2693 -823 -2659
rect -915 -2699 -823 -2693
rect -757 -2659 -665 -2653
rect -757 -2693 -728 -2659
rect -694 -2693 -665 -2659
rect -757 -2699 -665 -2693
rect -599 -2659 -507 -2653
rect -599 -2693 -570 -2659
rect -536 -2693 -507 -2659
rect -599 -2699 -507 -2693
rect -441 -2659 -349 -2653
rect -441 -2693 -412 -2659
rect -378 -2693 -349 -2659
rect -441 -2699 -349 -2693
rect -283 -2659 -191 -2653
rect -283 -2693 -254 -2659
rect -220 -2693 -191 -2659
rect -283 -2699 -191 -2693
rect -125 -2659 -33 -2653
rect -125 -2693 -96 -2659
rect -62 -2693 -33 -2659
rect -125 -2699 -33 -2693
rect 33 -2659 125 -2653
rect 33 -2693 62 -2659
rect 96 -2693 125 -2659
rect 33 -2699 125 -2693
rect 191 -2659 283 -2653
rect 191 -2693 220 -2659
rect 254 -2693 283 -2659
rect 191 -2699 283 -2693
rect 349 -2659 441 -2653
rect 349 -2693 378 -2659
rect 412 -2693 441 -2659
rect 349 -2699 441 -2693
rect 507 -2659 599 -2653
rect 507 -2693 536 -2659
rect 570 -2693 599 -2659
rect 507 -2699 599 -2693
rect 665 -2659 757 -2653
rect 665 -2693 694 -2659
rect 728 -2693 757 -2659
rect 665 -2699 757 -2693
rect 823 -2659 915 -2653
rect 823 -2693 852 -2659
rect 886 -2693 915 -2659
rect 823 -2699 915 -2693
rect 981 -2659 1073 -2653
rect 981 -2693 1010 -2659
rect 1044 -2693 1073 -2659
rect 981 -2699 1073 -2693
<< properties >>
string FIXED_BBOX -1220 -2778 1220 2778
<< end >>
