magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 24600 25950 24740 25990
rect 19760 21370 20200 21410
rect 24590 18790 24730 18830
rect 24590 17610 24730 17650
rect 19700 16820 20200 16860
rect 19750 15740 20210 15780
rect 19750 14940 20210 14980
rect 24590 10440 24730 10480
<< metal1 >>
rect 10240 22090 20210 22160
rect 20140 20480 20210 22090
rect 19740 19800 20080 19870
rect 20010 19200 20080 19800
rect 19990 19166 20100 19200
rect 19990 19114 20019 19166
rect 20071 19114 20100 19166
rect 19990 19080 20100 19114
rect 19700 19000 19910 19070
rect 19840 18650 19910 19000
rect 21660 18650 21770 18670
rect 19840 18641 21770 18650
rect 19840 18589 21689 18641
rect 21741 18589 21770 18641
rect 19840 18580 21770 18589
rect 21660 18560 21770 18580
rect 22120 18436 22230 18790
rect 22120 18384 22149 18436
rect 22201 18384 22230 18436
rect 22120 18360 22230 18384
rect 22820 18306 22930 18790
rect 26390 18750 26750 18800
rect 26650 18696 26750 18750
rect 26650 18644 26674 18696
rect 26726 18644 26750 18696
rect 26650 18620 26750 18644
rect 27350 18566 27450 18820
rect 27350 18514 27374 18566
rect 27426 18514 27450 18566
rect 27350 18490 27450 18514
rect 19750 17900 19820 18270
rect 22820 18254 22849 18306
rect 22901 18254 22930 18306
rect 22820 18230 22930 18254
rect 22120 18176 22230 18200
rect 22120 18124 22149 18176
rect 22201 18124 22230 18176
rect 21660 17900 21770 17920
rect 19750 17891 21770 17900
rect 19750 17839 21689 17891
rect 21741 17839 21770 17891
rect 19750 17830 21770 17839
rect 21660 17810 21770 17830
rect 22120 17610 22230 18124
rect 22820 18046 22930 18070
rect 22820 17994 22849 18046
rect 22901 17994 22930 18046
rect 22820 17610 22930 17994
rect 27350 17916 27450 17940
rect 27350 17864 27374 17916
rect 27426 17864 27450 17916
rect 26650 17786 26750 17810
rect 26650 17734 26674 17786
rect 26726 17734 26750 17786
rect 26650 17610 26750 17734
rect 27350 17610 27450 17864
rect 20130 17470 20240 17490
rect 19680 17461 20240 17470
rect 19680 17409 20159 17461
rect 20211 17409 20240 17461
rect 19680 17400 20240 17409
rect 20130 17380 20240 17400
rect 20140 13450 20202 15956
rect 10230 13380 20202 13450
<< via1 >>
rect 20019 19114 20071 19166
rect 21689 18589 21741 18641
rect 22149 18384 22201 18436
rect 26674 18644 26726 18696
rect 27374 18514 27426 18566
rect 22849 18254 22901 18306
rect 22149 18124 22201 18176
rect 21689 17839 21741 17891
rect 22849 17994 22901 18046
rect 27374 17864 27426 17916
rect 26674 17734 26726 17786
rect 20159 17409 20211 17461
<< metal2 >>
rect 18710 25420 20300 25860
rect 18710 20900 19000 25420
rect 20210 20923 20440 20930
rect 20210 20627 20217 20923
rect 20433 20627 20440 20923
rect 20210 20620 20440 20627
rect 19990 19168 20100 19200
rect 19990 19112 20017 19168
rect 20073 19112 20100 19168
rect 19990 19080 20100 19112
rect 22120 18696 29180 18720
rect 21660 18643 21770 18670
rect 21660 18587 21687 18643
rect 21743 18587 21770 18643
rect 22120 18644 26674 18696
rect 26726 18644 29180 18696
rect 22120 18620 29180 18644
rect 21660 18560 21770 18587
rect 22120 18566 29180 18590
rect 22120 18514 27374 18566
rect 27426 18514 29180 18566
rect 22120 18490 29180 18514
rect 22120 18436 29180 18460
rect 22120 18384 22149 18436
rect 22201 18384 29180 18436
rect 22120 18360 29180 18384
rect 22120 18306 29180 18330
rect 22120 18254 22849 18306
rect 22901 18254 29180 18306
rect 22120 18230 29180 18254
rect 22120 18176 29180 18200
rect 22120 18124 22149 18176
rect 22201 18124 29180 18176
rect 22120 18100 29180 18124
rect 22120 18046 29180 18070
rect 22120 17994 22849 18046
rect 22901 17994 29180 18046
rect 22120 17970 29180 17994
rect 21660 17893 21770 17920
rect 21660 17837 21687 17893
rect 21743 17837 21770 17893
rect 22120 17916 29180 17940
rect 22120 17864 27374 17916
rect 27426 17864 29180 17916
rect 22120 17840 29180 17864
rect 21660 17810 21770 17837
rect 22120 17786 29180 17810
rect 22120 17734 26674 17786
rect 26726 17734 29180 17786
rect 22120 17710 29180 17734
rect 20130 17463 20240 17490
rect 20130 17407 20157 17463
rect 20213 17407 20240 17463
rect 20130 17380 20240 17407
rect 17580 16983 19440 17020
rect 17580 16767 17632 16983
rect 17768 16767 19440 16983
rect 17580 16730 19440 16767
rect 10240 16000 19660 16430
rect 19230 15680 19660 16000
rect 17580 14378 18350 14420
rect 17580 14162 17642 14378
rect 17778 14162 18350 14378
rect 17580 14130 18350 14162
rect 19520 11010 19820 14420
rect 20650 13760 21050 15850
rect 20640 13470 21050 13760
rect 20640 13168 21040 13470
rect 20640 12872 20687 13168
rect 20983 12872 21040 13168
rect 20640 12820 21040 12872
rect 19520 10570 20250 11010
<< via2 >>
rect 20217 20627 20433 20923
rect 20017 19166 20073 19168
rect 20017 19114 20019 19166
rect 20019 19114 20071 19166
rect 20071 19114 20073 19166
rect 20017 19112 20073 19114
rect 21687 18641 21743 18643
rect 21687 18589 21689 18641
rect 21689 18589 21741 18641
rect 21741 18589 21743 18641
rect 21687 18587 21743 18589
rect 21687 17891 21743 17893
rect 21687 17839 21689 17891
rect 21689 17839 21741 17891
rect 21741 17839 21743 17891
rect 21687 17837 21743 17839
rect 20157 17461 20213 17463
rect 20157 17409 20159 17461
rect 20159 17409 20211 17461
rect 20211 17409 20213 17461
rect 20157 17407 20213 17409
rect 17632 16767 17768 16983
rect 17642 14162 17778 14378
rect 20687 12872 20983 13168
<< metal3 >>
rect 15670 20923 20500 20980
rect 15670 20627 20217 20923
rect 20433 20627 20500 20923
rect 15670 20580 20500 20627
rect 15670 20480 16440 20580
rect 15670 20270 16330 20480
rect 19990 19168 20410 19200
rect 19990 19112 20017 19168
rect 20073 19112 20410 19168
rect 19990 19080 20410 19112
rect 21150 18760 21450 26030
rect 22650 18670 22760 18830
rect 23350 18760 23650 26030
rect 21660 18643 22760 18670
rect 21660 18587 21687 18643
rect 21743 18587 22760 18643
rect 21660 18560 22760 18587
rect 25635 18330 25835 18939
rect 27680 18330 27880 18934
rect 19870 18100 27880 18330
rect 17540 16983 17840 17020
rect 17540 16767 17632 16983
rect 17768 16767 17840 16983
rect 10348 15604 10872 16712
rect 17540 14378 17840 16767
rect 17540 14162 17642 14378
rect 17778 14162 17840 14378
rect 17540 14130 17840 14162
rect 19870 13970 20070 18100
rect 21660 17893 22760 17920
rect 21660 17837 21687 17893
rect 21743 17837 22760 17893
rect 21660 17810 22760 17837
rect 20130 17463 20400 17490
rect 20130 17407 20157 17463
rect 20213 17407 20400 17463
rect 20130 17380 20400 17407
rect 19820 13570 20070 13970
rect 15850 13168 21040 13220
rect 15850 12872 20687 13168
rect 20983 12872 21040 13168
rect 15850 12820 21040 12872
rect 21150 10400 21450 17670
rect 22650 17570 22760 17810
rect 23350 10410 23650 17680
rect 25635 17490 25835 18100
rect 27680 17630 27880 18100
<< metal4 >>
rect 10225 20205 10250 20270
use buffer_amp  X1
timestamp 1663011646
transform 1 0 15140 0 1 17350
box 5000 1400 9520 8666
use buffer_amp  X2
timestamp 1663011646
transform 1 0 19660 0 -1 19081
box 5000 1400 9520 8666
use buffer_amp  X3
timestamp 1663011646
transform 1 0 15140 0 -1 19081
box 5000 1400 9520 8666
use buffer_amp  X4
timestamp 1663011646
transform 1 0 19660 0 1 17350
box 5000 1400 9520 8666
use amp_dec  X5
timestamp 1663011646
transform 0 1 9640 -1 0 26439
box 5000 590 10199 10186
use vop_dec  X6
timestamp 1663011646
transform 0 1 9830 -1 0 21409
box 5600 400 10899 9990
<< labels >>
rlabel metal2 s 10240 16000 19660 16430 4 VOP
port 1 nsew
rlabel metal3 s 15850 12820 20660 13220 4 GND
port 2 nsew
rlabel metal1 s 10230 13380 20140 13450 4 BIAS
port 3 nsew
rlabel metal3 s 21150 18760 21450 26030 4 OUT180
port 4 nsew
rlabel metal3 s 23350 18760 23650 26030 4 OUT0
port 5 nsew
rlabel metal3 s 21150 10400 21450 17670 4 OUT270
port 6 nsew
rlabel metal3 s 23350 10410 23650 17680 4 OUT90
port 7 nsew
rlabel locali s 19760 21370 20200 21410 4 SUB
port 8 nsew
rlabel metal1 s 10240 22090 20210 22160 4 BIAS
port 3 nsew
rlabel metal4 s 10225 20205 10250 20270 4 AMP
port 9 nsew
rlabel metal2 s 26730 18620 29180 18720 4 I4B
port 10 nsew
rlabel metal2 s 27430 18490 29180 18590 4 I4A
port 11 nsew
rlabel metal2 s 22210 18360 29180 18460 4 I1B
port 12 nsew
rlabel metal2 s 22910 18230 29180 18330 4 I1A
port 13 nsew
rlabel metal2 s 26740 18100 29180 18200 4 I3B
port 14 nsew
rlabel metal2 s 27440 17970 29180 18070 4 I3A
port 15 nsew
rlabel metal2 s 22920 17840 29180 17940 4 I2A
port 16 nsew
rlabel metal2 s 22220 17710 29180 17810 4 I2B
port 17 nsew
rlabel metal2 s 19520 10570 19820 14420 4 VDD
port 18 nsew
<< end >>
