magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -441 1712 441 1798
rect -441 -1712 -355 1712
rect 355 -1712 441 1712
rect -441 -1798 441 -1712
<< psubdiff >>
rect -415 1738 -289 1772
rect -255 1738 -221 1772
rect -187 1738 -153 1772
rect -119 1738 -85 1772
rect -51 1738 -17 1772
rect 17 1738 51 1772
rect 85 1738 119 1772
rect 153 1738 187 1772
rect 221 1738 255 1772
rect 289 1738 415 1772
rect -415 1649 -381 1738
rect 381 1649 415 1738
rect -415 1581 -381 1615
rect -415 1513 -381 1547
rect -415 1445 -381 1479
rect -415 1377 -381 1411
rect -415 1309 -381 1343
rect -415 1241 -381 1275
rect -415 1173 -381 1207
rect -415 1105 -381 1139
rect -415 1037 -381 1071
rect -415 969 -381 1003
rect -415 901 -381 935
rect -415 833 -381 867
rect -415 765 -381 799
rect -415 697 -381 731
rect -415 629 -381 663
rect -415 561 -381 595
rect -415 493 -381 527
rect -415 425 -381 459
rect -415 357 -381 391
rect -415 289 -381 323
rect -415 221 -381 255
rect -415 153 -381 187
rect -415 85 -381 119
rect -415 17 -381 51
rect -415 -51 -381 -17
rect -415 -119 -381 -85
rect -415 -187 -381 -153
rect -415 -255 -381 -221
rect -415 -323 -381 -289
rect -415 -391 -381 -357
rect -415 -459 -381 -425
rect -415 -527 -381 -493
rect -415 -595 -381 -561
rect -415 -663 -381 -629
rect -415 -731 -381 -697
rect -415 -799 -381 -765
rect -415 -867 -381 -833
rect -415 -935 -381 -901
rect -415 -1003 -381 -969
rect -415 -1071 -381 -1037
rect -415 -1139 -381 -1105
rect -415 -1207 -381 -1173
rect -415 -1275 -381 -1241
rect -415 -1343 -381 -1309
rect -415 -1411 -381 -1377
rect -415 -1479 -381 -1445
rect -415 -1547 -381 -1513
rect -415 -1615 -381 -1581
rect 381 1581 415 1615
rect 381 1513 415 1547
rect 381 1445 415 1479
rect 381 1377 415 1411
rect 381 1309 415 1343
rect 381 1241 415 1275
rect 381 1173 415 1207
rect 381 1105 415 1139
rect 381 1037 415 1071
rect 381 969 415 1003
rect 381 901 415 935
rect 381 833 415 867
rect 381 765 415 799
rect 381 697 415 731
rect 381 629 415 663
rect 381 561 415 595
rect 381 493 415 527
rect 381 425 415 459
rect 381 357 415 391
rect 381 289 415 323
rect 381 221 415 255
rect 381 153 415 187
rect 381 85 415 119
rect 381 17 415 51
rect 381 -51 415 -17
rect 381 -119 415 -85
rect 381 -187 415 -153
rect 381 -255 415 -221
rect 381 -323 415 -289
rect 381 -391 415 -357
rect 381 -459 415 -425
rect 381 -527 415 -493
rect 381 -595 415 -561
rect 381 -663 415 -629
rect 381 -731 415 -697
rect 381 -799 415 -765
rect 381 -867 415 -833
rect 381 -935 415 -901
rect 381 -1003 415 -969
rect 381 -1071 415 -1037
rect 381 -1139 415 -1105
rect 381 -1207 415 -1173
rect 381 -1275 415 -1241
rect 381 -1343 415 -1309
rect 381 -1411 415 -1377
rect 381 -1479 415 -1445
rect 381 -1547 415 -1513
rect 381 -1615 415 -1581
rect -415 -1738 -381 -1649
rect 381 -1738 415 -1649
rect -415 -1772 -289 -1738
rect -255 -1772 -221 -1738
rect -187 -1772 -153 -1738
rect -119 -1772 -85 -1738
rect -51 -1772 -17 -1738
rect 17 -1772 51 -1738
rect 85 -1772 119 -1738
rect 153 -1772 187 -1738
rect 221 -1772 255 -1738
rect 289 -1772 415 -1738
<< psubdiffcont >>
rect -289 1738 -255 1772
rect -221 1738 -187 1772
rect -153 1738 -119 1772
rect -85 1738 -51 1772
rect -17 1738 17 1772
rect 51 1738 85 1772
rect 119 1738 153 1772
rect 187 1738 221 1772
rect 255 1738 289 1772
rect -415 1615 -381 1649
rect -415 1547 -381 1581
rect -415 1479 -381 1513
rect -415 1411 -381 1445
rect -415 1343 -381 1377
rect -415 1275 -381 1309
rect -415 1207 -381 1241
rect -415 1139 -381 1173
rect -415 1071 -381 1105
rect -415 1003 -381 1037
rect -415 935 -381 969
rect -415 867 -381 901
rect -415 799 -381 833
rect -415 731 -381 765
rect -415 663 -381 697
rect -415 595 -381 629
rect -415 527 -381 561
rect -415 459 -381 493
rect -415 391 -381 425
rect -415 323 -381 357
rect -415 255 -381 289
rect -415 187 -381 221
rect -415 119 -381 153
rect -415 51 -381 85
rect -415 -17 -381 17
rect -415 -85 -381 -51
rect -415 -153 -381 -119
rect -415 -221 -381 -187
rect -415 -289 -381 -255
rect -415 -357 -381 -323
rect -415 -425 -381 -391
rect -415 -493 -381 -459
rect -415 -561 -381 -527
rect -415 -629 -381 -595
rect -415 -697 -381 -663
rect -415 -765 -381 -731
rect -415 -833 -381 -799
rect -415 -901 -381 -867
rect -415 -969 -381 -935
rect -415 -1037 -381 -1003
rect -415 -1105 -381 -1071
rect -415 -1173 -381 -1139
rect -415 -1241 -381 -1207
rect -415 -1309 -381 -1275
rect -415 -1377 -381 -1343
rect -415 -1445 -381 -1411
rect -415 -1513 -381 -1479
rect -415 -1581 -381 -1547
rect -415 -1649 -381 -1615
rect 381 1615 415 1649
rect 381 1547 415 1581
rect 381 1479 415 1513
rect 381 1411 415 1445
rect 381 1343 415 1377
rect 381 1275 415 1309
rect 381 1207 415 1241
rect 381 1139 415 1173
rect 381 1071 415 1105
rect 381 1003 415 1037
rect 381 935 415 969
rect 381 867 415 901
rect 381 799 415 833
rect 381 731 415 765
rect 381 663 415 697
rect 381 595 415 629
rect 381 527 415 561
rect 381 459 415 493
rect 381 391 415 425
rect 381 323 415 357
rect 381 255 415 289
rect 381 187 415 221
rect 381 119 415 153
rect 381 51 415 85
rect 381 -17 415 17
rect 381 -85 415 -51
rect 381 -153 415 -119
rect 381 -221 415 -187
rect 381 -289 415 -255
rect 381 -357 415 -323
rect 381 -425 415 -391
rect 381 -493 415 -459
rect 381 -561 415 -527
rect 381 -629 415 -595
rect 381 -697 415 -663
rect 381 -765 415 -731
rect 381 -833 415 -799
rect 381 -901 415 -867
rect 381 -969 415 -935
rect 381 -1037 415 -1003
rect 381 -1105 415 -1071
rect 381 -1173 415 -1139
rect 381 -1241 415 -1207
rect 381 -1309 415 -1275
rect 381 -1377 415 -1343
rect 381 -1445 415 -1411
rect 381 -1513 415 -1479
rect 381 -1581 415 -1547
rect 381 -1649 415 -1615
rect -289 -1772 -255 -1738
rect -221 -1772 -187 -1738
rect -153 -1772 -119 -1738
rect -85 -1772 -51 -1738
rect -17 -1772 17 -1738
rect 51 -1772 85 -1738
rect 119 -1772 153 -1738
rect 187 -1772 221 -1738
rect 255 -1772 289 -1738
<< xpolycontact >>
rect -285 1210 285 1642
rect -285 -1642 285 -1210
<< ppolyres >>
rect -285 -1210 285 1210
<< locali >>
rect -415 1738 -289 1772
rect -255 1738 -221 1772
rect -187 1738 -153 1772
rect -119 1738 -85 1772
rect -51 1738 -17 1772
rect 17 1738 51 1772
rect 85 1738 119 1772
rect 153 1738 187 1772
rect 221 1738 255 1772
rect 289 1738 415 1772
rect -415 1649 -381 1738
rect 381 1649 415 1738
rect -415 1581 -381 1615
rect -415 1513 -381 1547
rect -415 1445 -381 1479
rect -415 1377 -381 1411
rect -415 1309 -381 1343
rect -415 1241 -381 1275
rect 381 1581 415 1615
rect 381 1513 415 1547
rect 381 1445 415 1479
rect 381 1377 415 1411
rect 381 1309 415 1343
rect 381 1241 415 1275
rect -415 1173 -381 1207
rect -415 1105 -381 1139
rect -415 1037 -381 1071
rect -415 969 -381 1003
rect -415 901 -381 935
rect -415 833 -381 867
rect -415 765 -381 799
rect -415 697 -381 731
rect -415 629 -381 663
rect -415 561 -381 595
rect -415 493 -381 527
rect -415 425 -381 459
rect -415 357 -381 391
rect -415 289 -381 323
rect -415 221 -381 255
rect -415 153 -381 187
rect -415 85 -381 119
rect -415 17 -381 51
rect -415 -51 -381 -17
rect -415 -119 -381 -85
rect -415 -187 -381 -153
rect -415 -255 -381 -221
rect -415 -323 -381 -289
rect -415 -391 -381 -357
rect -415 -459 -381 -425
rect -415 -527 -381 -493
rect -415 -595 -381 -561
rect -415 -663 -381 -629
rect -415 -731 -381 -697
rect -415 -799 -381 -765
rect -415 -867 -381 -833
rect -415 -935 -381 -901
rect -415 -1003 -381 -969
rect -415 -1071 -381 -1037
rect -415 -1139 -381 -1105
rect -415 -1207 -381 -1173
rect 381 1173 415 1207
rect 381 1105 415 1139
rect 381 1037 415 1071
rect 381 969 415 1003
rect 381 901 415 935
rect 381 833 415 867
rect 381 765 415 799
rect 381 697 415 731
rect 381 629 415 663
rect 381 561 415 595
rect 381 493 415 527
rect 381 425 415 459
rect 381 357 415 391
rect 381 289 415 323
rect 381 221 415 255
rect 381 153 415 187
rect 381 85 415 119
rect 381 17 415 51
rect 381 -51 415 -17
rect 381 -119 415 -85
rect 381 -187 415 -153
rect 381 -255 415 -221
rect 381 -323 415 -289
rect 381 -391 415 -357
rect 381 -459 415 -425
rect 381 -527 415 -493
rect 381 -595 415 -561
rect 381 -663 415 -629
rect 381 -731 415 -697
rect 381 -799 415 -765
rect 381 -867 415 -833
rect 381 -935 415 -901
rect 381 -1003 415 -969
rect 381 -1071 415 -1037
rect 381 -1139 415 -1105
rect 381 -1207 415 -1173
rect -415 -1275 -381 -1241
rect -415 -1343 -381 -1309
rect -415 -1411 -381 -1377
rect -415 -1479 -381 -1445
rect -415 -1547 -381 -1513
rect -415 -1615 -381 -1581
rect 381 -1275 415 -1241
rect 381 -1343 415 -1309
rect 381 -1411 415 -1377
rect 381 -1479 415 -1445
rect 381 -1547 415 -1513
rect 381 -1615 415 -1581
rect -415 -1738 -381 -1649
rect 381 -1738 415 -1649
rect -415 -1772 -289 -1738
rect -255 -1772 -221 -1738
rect -187 -1772 -153 -1738
rect -119 -1772 -85 -1738
rect -51 -1772 -17 -1738
rect 17 -1772 51 -1738
rect 85 -1772 119 -1738
rect 153 -1772 187 -1738
rect 221 -1772 255 -1738
rect 289 -1772 415 -1738
<< viali >>
rect -269 1228 269 1622
rect -269 -1623 269 -1229
<< metal1 >>
rect -281 1622 281 1630
rect -281 1228 -269 1622
rect 269 1228 281 1622
rect -281 1221 281 1228
rect -281 -1229 281 -1221
rect -281 -1623 -269 -1229
rect 269 -1623 281 -1229
rect -281 -1630 281 -1623
<< properties >>
string FIXED_BBOX -398 -1755 398 1755
<< end >>
