magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -729 2142 729 2228
rect -729 -2142 -643 2142
rect 643 -2142 729 2142
rect -729 -2228 729 -2142
<< psubdiff >>
rect -703 2168 -595 2202
rect -561 2168 -527 2202
rect -493 2168 -459 2202
rect -425 2168 -391 2202
rect -357 2168 -323 2202
rect -289 2168 -255 2202
rect -221 2168 -187 2202
rect -153 2168 -119 2202
rect -85 2168 -51 2202
rect -17 2168 17 2202
rect 51 2168 85 2202
rect 119 2168 153 2202
rect 187 2168 221 2202
rect 255 2168 289 2202
rect 323 2168 357 2202
rect 391 2168 425 2202
rect 459 2168 493 2202
rect 527 2168 561 2202
rect 595 2168 703 2202
rect -703 2091 -669 2168
rect 669 2091 703 2168
rect -703 2023 -669 2057
rect -703 1955 -669 1989
rect -703 1887 -669 1921
rect -703 1819 -669 1853
rect -703 1751 -669 1785
rect -703 1683 -669 1717
rect -703 1615 -669 1649
rect -703 1547 -669 1581
rect -703 1479 -669 1513
rect -703 1411 -669 1445
rect -703 1343 -669 1377
rect -703 1275 -669 1309
rect -703 1207 -669 1241
rect -703 1139 -669 1173
rect -703 1071 -669 1105
rect -703 1003 -669 1037
rect -703 935 -669 969
rect -703 867 -669 901
rect -703 799 -669 833
rect -703 731 -669 765
rect -703 663 -669 697
rect -703 595 -669 629
rect -703 527 -669 561
rect -703 459 -669 493
rect -703 391 -669 425
rect -703 323 -669 357
rect -703 255 -669 289
rect -703 187 -669 221
rect -703 119 -669 153
rect -703 51 -669 85
rect -703 -17 -669 17
rect -703 -85 -669 -51
rect -703 -153 -669 -119
rect -703 -221 -669 -187
rect -703 -289 -669 -255
rect -703 -357 -669 -323
rect -703 -425 -669 -391
rect -703 -493 -669 -459
rect -703 -561 -669 -527
rect -703 -629 -669 -595
rect -703 -697 -669 -663
rect -703 -765 -669 -731
rect -703 -833 -669 -799
rect -703 -901 -669 -867
rect -703 -969 -669 -935
rect -703 -1037 -669 -1003
rect -703 -1105 -669 -1071
rect -703 -1173 -669 -1139
rect -703 -1241 -669 -1207
rect -703 -1309 -669 -1275
rect -703 -1377 -669 -1343
rect -703 -1445 -669 -1411
rect -703 -1513 -669 -1479
rect -703 -1581 -669 -1547
rect -703 -1649 -669 -1615
rect -703 -1717 -669 -1683
rect -703 -1785 -669 -1751
rect -703 -1853 -669 -1819
rect -703 -1921 -669 -1887
rect -703 -1989 -669 -1955
rect -703 -2057 -669 -2023
rect 669 2023 703 2057
rect 669 1955 703 1989
rect 669 1887 703 1921
rect 669 1819 703 1853
rect 669 1751 703 1785
rect 669 1683 703 1717
rect 669 1615 703 1649
rect 669 1547 703 1581
rect 669 1479 703 1513
rect 669 1411 703 1445
rect 669 1343 703 1377
rect 669 1275 703 1309
rect 669 1207 703 1241
rect 669 1139 703 1173
rect 669 1071 703 1105
rect 669 1003 703 1037
rect 669 935 703 969
rect 669 867 703 901
rect 669 799 703 833
rect 669 731 703 765
rect 669 663 703 697
rect 669 595 703 629
rect 669 527 703 561
rect 669 459 703 493
rect 669 391 703 425
rect 669 323 703 357
rect 669 255 703 289
rect 669 187 703 221
rect 669 119 703 153
rect 669 51 703 85
rect 669 -17 703 17
rect 669 -85 703 -51
rect 669 -153 703 -119
rect 669 -221 703 -187
rect 669 -289 703 -255
rect 669 -357 703 -323
rect 669 -425 703 -391
rect 669 -493 703 -459
rect 669 -561 703 -527
rect 669 -629 703 -595
rect 669 -697 703 -663
rect 669 -765 703 -731
rect 669 -833 703 -799
rect 669 -901 703 -867
rect 669 -969 703 -935
rect 669 -1037 703 -1003
rect 669 -1105 703 -1071
rect 669 -1173 703 -1139
rect 669 -1241 703 -1207
rect 669 -1309 703 -1275
rect 669 -1377 703 -1343
rect 669 -1445 703 -1411
rect 669 -1513 703 -1479
rect 669 -1581 703 -1547
rect 669 -1649 703 -1615
rect 669 -1717 703 -1683
rect 669 -1785 703 -1751
rect 669 -1853 703 -1819
rect 669 -1921 703 -1887
rect 669 -1989 703 -1955
rect 669 -2057 703 -2023
rect -703 -2168 -669 -2091
rect 669 -2168 703 -2091
rect -703 -2202 -595 -2168
rect -561 -2202 -527 -2168
rect -493 -2202 -459 -2168
rect -425 -2202 -391 -2168
rect -357 -2202 -323 -2168
rect -289 -2202 -255 -2168
rect -221 -2202 -187 -2168
rect -153 -2202 -119 -2168
rect -85 -2202 -51 -2168
rect -17 -2202 17 -2168
rect 51 -2202 85 -2168
rect 119 -2202 153 -2168
rect 187 -2202 221 -2168
rect 255 -2202 289 -2168
rect 323 -2202 357 -2168
rect 391 -2202 425 -2168
rect 459 -2202 493 -2168
rect 527 -2202 561 -2168
rect 595 -2202 703 -2168
<< psubdiffcont >>
rect -595 2168 -561 2202
rect -527 2168 -493 2202
rect -459 2168 -425 2202
rect -391 2168 -357 2202
rect -323 2168 -289 2202
rect -255 2168 -221 2202
rect -187 2168 -153 2202
rect -119 2168 -85 2202
rect -51 2168 -17 2202
rect 17 2168 51 2202
rect 85 2168 119 2202
rect 153 2168 187 2202
rect 221 2168 255 2202
rect 289 2168 323 2202
rect 357 2168 391 2202
rect 425 2168 459 2202
rect 493 2168 527 2202
rect 561 2168 595 2202
rect -703 2057 -669 2091
rect -703 1989 -669 2023
rect -703 1921 -669 1955
rect -703 1853 -669 1887
rect -703 1785 -669 1819
rect -703 1717 -669 1751
rect -703 1649 -669 1683
rect -703 1581 -669 1615
rect -703 1513 -669 1547
rect -703 1445 -669 1479
rect -703 1377 -669 1411
rect -703 1309 -669 1343
rect -703 1241 -669 1275
rect -703 1173 -669 1207
rect -703 1105 -669 1139
rect -703 1037 -669 1071
rect -703 969 -669 1003
rect -703 901 -669 935
rect -703 833 -669 867
rect -703 765 -669 799
rect -703 697 -669 731
rect -703 629 -669 663
rect -703 561 -669 595
rect -703 493 -669 527
rect -703 425 -669 459
rect -703 357 -669 391
rect -703 289 -669 323
rect -703 221 -669 255
rect -703 153 -669 187
rect -703 85 -669 119
rect -703 17 -669 51
rect -703 -51 -669 -17
rect -703 -119 -669 -85
rect -703 -187 -669 -153
rect -703 -255 -669 -221
rect -703 -323 -669 -289
rect -703 -391 -669 -357
rect -703 -459 -669 -425
rect -703 -527 -669 -493
rect -703 -595 -669 -561
rect -703 -663 -669 -629
rect -703 -731 -669 -697
rect -703 -799 -669 -765
rect -703 -867 -669 -833
rect -703 -935 -669 -901
rect -703 -1003 -669 -969
rect -703 -1071 -669 -1037
rect -703 -1139 -669 -1105
rect -703 -1207 -669 -1173
rect -703 -1275 -669 -1241
rect -703 -1343 -669 -1309
rect -703 -1411 -669 -1377
rect -703 -1479 -669 -1445
rect -703 -1547 -669 -1513
rect -703 -1615 -669 -1581
rect -703 -1683 -669 -1649
rect -703 -1751 -669 -1717
rect -703 -1819 -669 -1785
rect -703 -1887 -669 -1853
rect -703 -1955 -669 -1921
rect -703 -2023 -669 -1989
rect -703 -2091 -669 -2057
rect 669 2057 703 2091
rect 669 1989 703 2023
rect 669 1921 703 1955
rect 669 1853 703 1887
rect 669 1785 703 1819
rect 669 1717 703 1751
rect 669 1649 703 1683
rect 669 1581 703 1615
rect 669 1513 703 1547
rect 669 1445 703 1479
rect 669 1377 703 1411
rect 669 1309 703 1343
rect 669 1241 703 1275
rect 669 1173 703 1207
rect 669 1105 703 1139
rect 669 1037 703 1071
rect 669 969 703 1003
rect 669 901 703 935
rect 669 833 703 867
rect 669 765 703 799
rect 669 697 703 731
rect 669 629 703 663
rect 669 561 703 595
rect 669 493 703 527
rect 669 425 703 459
rect 669 357 703 391
rect 669 289 703 323
rect 669 221 703 255
rect 669 153 703 187
rect 669 85 703 119
rect 669 17 703 51
rect 669 -51 703 -17
rect 669 -119 703 -85
rect 669 -187 703 -153
rect 669 -255 703 -221
rect 669 -323 703 -289
rect 669 -391 703 -357
rect 669 -459 703 -425
rect 669 -527 703 -493
rect 669 -595 703 -561
rect 669 -663 703 -629
rect 669 -731 703 -697
rect 669 -799 703 -765
rect 669 -867 703 -833
rect 669 -935 703 -901
rect 669 -1003 703 -969
rect 669 -1071 703 -1037
rect 669 -1139 703 -1105
rect 669 -1207 703 -1173
rect 669 -1275 703 -1241
rect 669 -1343 703 -1309
rect 669 -1411 703 -1377
rect 669 -1479 703 -1445
rect 669 -1547 703 -1513
rect 669 -1615 703 -1581
rect 669 -1683 703 -1649
rect 669 -1751 703 -1717
rect 669 -1819 703 -1785
rect 669 -1887 703 -1853
rect 669 -1955 703 -1921
rect 669 -2023 703 -1989
rect 669 -2091 703 -2057
rect -595 -2202 -561 -2168
rect -527 -2202 -493 -2168
rect -459 -2202 -425 -2168
rect -391 -2202 -357 -2168
rect -323 -2202 -289 -2168
rect -255 -2202 -221 -2168
rect -187 -2202 -153 -2168
rect -119 -2202 -85 -2168
rect -51 -2202 -17 -2168
rect 17 -2202 51 -2168
rect 85 -2202 119 -2168
rect 153 -2202 187 -2168
rect 221 -2202 255 -2168
rect 289 -2202 323 -2168
rect 357 -2202 391 -2168
rect 425 -2202 459 -2168
rect 493 -2202 527 -2168
rect 561 -2202 595 -2168
<< xpolycontact >>
rect -573 1640 573 2072
rect -573 -2072 573 -1640
<< ppolyres >>
rect -573 -1640 573 1640
<< locali >>
rect -703 2168 -595 2202
rect -561 2168 -527 2202
rect -493 2168 -459 2202
rect -425 2168 -391 2202
rect -357 2168 -323 2202
rect -289 2168 -255 2202
rect -221 2168 -187 2202
rect -153 2168 -119 2202
rect -85 2168 -51 2202
rect -17 2168 17 2202
rect 51 2168 85 2202
rect 119 2168 153 2202
rect 187 2168 221 2202
rect 255 2168 289 2202
rect 323 2168 357 2202
rect 391 2168 425 2202
rect 459 2168 493 2202
rect 527 2168 561 2202
rect 595 2168 703 2202
rect -703 2091 -669 2168
rect 669 2091 703 2168
rect -703 2023 -669 2057
rect -703 1955 -669 1989
rect -703 1887 -669 1921
rect -703 1819 -669 1853
rect -703 1751 -669 1785
rect -703 1683 -669 1717
rect -703 1615 -669 1649
rect 669 2023 703 2057
rect 669 1955 703 1989
rect 669 1887 703 1921
rect 669 1819 703 1853
rect 669 1751 703 1785
rect 669 1683 703 1717
rect -703 1547 -669 1581
rect -703 1479 -669 1513
rect -703 1411 -669 1445
rect -703 1343 -669 1377
rect -703 1275 -669 1309
rect -703 1207 -669 1241
rect -703 1139 -669 1173
rect -703 1071 -669 1105
rect -703 1003 -669 1037
rect -703 935 -669 969
rect -703 867 -669 901
rect -703 799 -669 833
rect -703 731 -669 765
rect -703 663 -669 697
rect -703 595 -669 629
rect -703 527 -669 561
rect -703 459 -669 493
rect -703 391 -669 425
rect -703 323 -669 357
rect -703 255 -669 289
rect -703 187 -669 221
rect -703 119 -669 153
rect -703 51 -669 85
rect -703 -17 -669 17
rect -703 -85 -669 -51
rect -703 -153 -669 -119
rect -703 -221 -669 -187
rect -703 -289 -669 -255
rect -703 -357 -669 -323
rect -703 -425 -669 -391
rect -703 -493 -669 -459
rect -703 -561 -669 -527
rect -703 -629 -669 -595
rect -703 -697 -669 -663
rect -703 -765 -669 -731
rect -703 -833 -669 -799
rect -703 -901 -669 -867
rect -703 -969 -669 -935
rect -703 -1037 -669 -1003
rect -703 -1105 -669 -1071
rect -703 -1173 -669 -1139
rect -703 -1241 -669 -1207
rect -703 -1309 -669 -1275
rect -703 -1377 -669 -1343
rect -703 -1445 -669 -1411
rect -703 -1513 -669 -1479
rect -703 -1581 -669 -1547
rect -703 -1649 -669 -1615
rect 669 1615 703 1649
rect 669 1547 703 1581
rect 669 1479 703 1513
rect 669 1411 703 1445
rect 669 1343 703 1377
rect 669 1275 703 1309
rect 669 1207 703 1241
rect 669 1139 703 1173
rect 669 1071 703 1105
rect 669 1003 703 1037
rect 669 935 703 969
rect 669 867 703 901
rect 669 799 703 833
rect 669 731 703 765
rect 669 663 703 697
rect 669 595 703 629
rect 669 527 703 561
rect 669 459 703 493
rect 669 391 703 425
rect 669 323 703 357
rect 669 255 703 289
rect 669 187 703 221
rect 669 119 703 153
rect 669 51 703 85
rect 669 -17 703 17
rect 669 -85 703 -51
rect 669 -153 703 -119
rect 669 -221 703 -187
rect 669 -289 703 -255
rect 669 -357 703 -323
rect 669 -425 703 -391
rect 669 -493 703 -459
rect 669 -561 703 -527
rect 669 -629 703 -595
rect 669 -697 703 -663
rect 669 -765 703 -731
rect 669 -833 703 -799
rect 669 -901 703 -867
rect 669 -969 703 -935
rect 669 -1037 703 -1003
rect 669 -1105 703 -1071
rect 669 -1173 703 -1139
rect 669 -1241 703 -1207
rect 669 -1309 703 -1275
rect 669 -1377 703 -1343
rect 669 -1445 703 -1411
rect 669 -1513 703 -1479
rect 669 -1581 703 -1547
rect -703 -1717 -669 -1683
rect -703 -1785 -669 -1751
rect -703 -1853 -669 -1819
rect -703 -1921 -669 -1887
rect -703 -1989 -669 -1955
rect -703 -2057 -669 -2023
rect 669 -1649 703 -1615
rect 669 -1717 703 -1683
rect 669 -1785 703 -1751
rect 669 -1853 703 -1819
rect 669 -1921 703 -1887
rect 669 -1989 703 -1955
rect 669 -2057 703 -2023
rect -703 -2168 -669 -2091
rect 669 -2168 703 -2091
rect -703 -2202 -595 -2168
rect -561 -2202 -527 -2168
rect -493 -2202 -459 -2168
rect -425 -2202 -391 -2168
rect -357 -2202 -323 -2168
rect -289 -2202 -255 -2168
rect -221 -2202 -187 -2168
rect -153 -2202 -119 -2168
rect -85 -2202 -51 -2168
rect -17 -2202 17 -2168
rect 51 -2202 85 -2168
rect 119 -2202 153 -2168
rect 187 -2202 221 -2168
rect 255 -2202 289 -2168
rect 323 -2202 357 -2168
rect 391 -2202 425 -2168
rect 459 -2202 493 -2168
rect 527 -2202 561 -2168
rect 595 -2202 703 -2168
<< viali >>
rect -557 1658 557 2052
rect -557 -2053 557 -1659
<< metal1 >>
rect -569 2052 569 2060
rect -569 1658 -557 2052
rect 557 1658 569 2052
rect -569 1651 569 1658
rect -569 -1659 569 -1651
rect -569 -2053 -557 -1659
rect 557 -2053 569 -1659
rect -569 -2060 569 -2053
<< properties >>
string FIXED_BBOX -686 -2185 686 2185
<< end >>
