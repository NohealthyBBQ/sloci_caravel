magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 12290 11270 12670 11305
rect 12290 8660 12670 8695
rect 10175 7140 10215 8395
rect 11345 7140 11385 8395
rect 13575 7140 13615 8395
rect 14750 7140 14790 8395
rect 12290 6840 12670 6875
rect 12290 4230 12670 4265
<< metal2 >>
rect 12280 12036 14415 12111
rect 15735 12035 16085 12110
rect 15910 11823 15990 11835
rect 15910 11767 15922 11823
rect 15978 11767 15990 11823
rect 15910 11750 15990 11767
rect 15810 11458 15890 11470
rect 15810 11402 15822 11458
rect 15878 11402 15890 11458
rect 15810 11390 15890 11402
rect 9185 8253 10505 8275
rect 9185 8197 10432 8253
rect 10488 8197 10505 8253
rect 9185 8175 10505 8197
rect 10575 8145 10675 8330
rect 11130 8275 11230 8325
rect 13625 8320 13630 8380
rect 13635 8373 13695 8375
rect 13635 8320 13637 8373
rect 13625 8317 13637 8320
rect 13693 8320 13695 8373
rect 14660 8368 14740 8395
rect 13693 8317 13705 8320
rect 13625 8305 13705 8317
rect 14660 8312 14672 8368
rect 14728 8312 14740 8368
rect 14660 8305 14740 8312
rect 10765 8253 15760 8275
rect 10765 8197 10782 8253
rect 10838 8197 12792 8253
rect 12848 8197 15760 8253
rect 10765 8175 15760 8197
rect 9185 8125 15760 8145
rect 9185 8069 14862 8125
rect 14918 8069 15760 8125
rect 9185 8045 15760 8069
rect 9185 7993 15760 8015
rect 9185 7937 10237 7993
rect 10293 7937 15760 7993
rect 9185 7915 15760 7937
rect 9185 7863 15760 7885
rect 9185 7807 11272 7863
rect 11328 7807 15760 7863
rect 9185 7785 15760 7807
rect 9185 7733 15760 7755
rect 9185 7677 13637 7733
rect 13693 7677 15760 7733
rect 9185 7655 15760 7677
rect 9185 7603 15760 7625
rect 9185 7547 14672 7603
rect 14728 7547 15760 7603
rect 9185 7525 15760 7547
rect 9180 7473 15760 7495
rect 9180 7417 12117 7473
rect 12173 7417 15760 7473
rect 9180 7395 15760 7417
rect 9175 7343 14190 7365
rect 9175 7287 9857 7343
rect 9913 7287 14122 7343
rect 14178 7287 14190 7343
rect 9175 7265 14190 7287
rect 10225 7223 10305 7235
rect 10225 7167 10237 7223
rect 10293 7167 10305 7223
rect 10225 7140 10305 7167
rect 11260 7223 11340 7235
rect 11260 7167 11272 7223
rect 11328 7167 11340 7223
rect 13755 7210 13830 7265
rect 14285 7215 14360 7395
rect 14460 7343 15760 7365
rect 14460 7287 14472 7343
rect 14528 7287 15760 7343
rect 14460 7265 15760 7287
rect 11260 7155 11340 7167
rect 15825 4173 15890 11390
rect 15825 4145 15827 4173
rect 15815 4117 15827 4145
rect 15883 4117 15890 4173
rect 15815 4105 15890 4117
rect 15925 3770 15990 11750
rect 15910 3758 15990 3770
rect 15910 3702 15922 3758
rect 15978 3702 15990 3758
rect 15910 3685 15990 3702
rect 16020 3500 16085 12035
rect 12350 3425 13635 3500
rect 15730 3425 16085 3500
<< via2 >>
rect 15922 11767 15978 11823
rect 15822 11402 15878 11458
rect 10432 8197 10488 8253
rect 13637 8317 13693 8373
rect 14672 8312 14728 8368
rect 10782 8197 10838 8253
rect 12792 8197 12848 8253
rect 14862 8069 14918 8125
rect 10237 7937 10293 7993
rect 11272 7807 11328 7863
rect 13637 7677 13693 7733
rect 14672 7547 14728 7603
rect 12117 7417 12173 7473
rect 9857 7287 9913 7343
rect 14122 7287 14178 7343
rect 10237 7167 10293 7223
rect 11272 7167 11328 7223
rect 14472 7287 14528 7343
rect 15827 4117 15883 4173
rect 15922 3702 15978 3758
<< metal3 >>
rect 12355 11705 12775 12005
rect 15735 11823 15990 11835
rect 15735 11775 15922 11823
rect 15910 11767 15922 11775
rect 15978 11767 15990 11823
rect 15910 11750 15990 11767
rect 12350 11295 13540 11595
rect 15710 11458 15890 11470
rect 15710 11402 15822 11458
rect 15878 11402 15890 11458
rect 15710 11390 15890 11402
rect 10225 7993 10305 8460
rect 10415 8253 10855 8275
rect 10415 8197 10432 8253
rect 10488 8197 10782 8253
rect 10838 8197 10855 8253
rect 10415 8175 10855 8197
rect 10225 7937 10237 7993
rect 10293 7937 10305 7993
rect 9835 7343 9935 7365
rect 9835 7287 9857 7343
rect 9913 7287 9935 7343
rect 9835 6790 9935 7287
rect 10225 7223 10305 7937
rect 10225 7167 10237 7223
rect 10293 7167 10305 7223
rect 10225 7155 10305 7167
rect 11260 7863 11340 8445
rect 12770 8253 12870 8780
rect 12770 8197 12792 8253
rect 12848 8197 12870 8253
rect 12770 8175 12870 8197
rect 13625 8373 13705 8380
rect 13625 8317 13637 8373
rect 13693 8317 13705 8373
rect 11260 7807 11272 7863
rect 11328 7807 11340 7863
rect 11260 7223 11340 7807
rect 13625 7733 13705 8317
rect 13625 7677 13637 7733
rect 13693 7677 13705 7733
rect 11260 7167 11272 7223
rect 11328 7167 11340 7223
rect 11260 7155 11340 7167
rect 12095 7473 12195 7495
rect 12095 7417 12117 7473
rect 12173 7417 12195 7473
rect 12095 6790 12195 7417
rect 13625 7065 13705 7677
rect 14660 8368 14740 8380
rect 14660 8312 14672 8368
rect 14728 8312 14740 8368
rect 14660 7603 14740 8312
rect 14840 8125 14940 8740
rect 14840 8069 14862 8125
rect 14918 8069 14940 8125
rect 14840 8045 14940 8069
rect 14660 7547 14672 7603
rect 14728 7547 14740 7603
rect 14110 7343 14540 7365
rect 14110 7287 14122 7343
rect 14178 7287 14472 7343
rect 14528 7287 14540 7343
rect 14110 7265 14540 7287
rect 14660 7085 14740 7547
rect 12355 4075 13525 4240
rect 15725 4173 15890 4180
rect 15725 4120 15827 4173
rect 15750 4117 15827 4120
rect 15883 4117 15890 4173
rect 15750 4105 15890 4117
rect 12355 3940 13525 4005
rect 12355 3810 13525 3830
rect 12355 3550 12787 3810
rect 13317 3550 13525 3810
rect 15910 3758 15990 3770
rect 15910 3755 15922 3758
rect 15695 3702 15922 3755
rect 15978 3702 15990 3758
rect 15695 3685 15990 3702
rect 12355 3530 13525 3550
use core_osc_amp  X1
timestamp 1663011646
transform -1 0 14762 0 -1 12340
box 2400 230 5552 4020
use core_osc_amp  X2
timestamp 1663011646
transform -1 0 14762 0 1 3195
box 2400 230 5552 4020
use core_osc_amp  X3
timestamp 1663011646
transform -1 0 18162 0 1 3195
box 2400 230 5552 4020
use core_osc_amp  X4
timestamp 1663011646
transform -1 0 18162 0 -1 12340
box 2400 230 5552 4020
<< labels >>
rlabel metal2 s 9185 8045 14850 8145 4 S4A
port 1 nsew
rlabel metal2 s 9185 7915 10235 8015 4 S1B
port 2 nsew
rlabel metal2 s 9185 7785 11270 7885 4 S1A
port 3 nsew
rlabel metal2 s 9185 7655 13635 7755 4 S3B
port 4 nsew
rlabel metal2 s 9185 7525 14670 7625 4 S3A
port 5 nsew
rlabel metal2 s 9180 7395 12100 7495 4 S2A
port 6 nsew
rlabel metal2 s 9175 7265 9845 7365 4 S2B
port 7 nsew
rlabel metal2 s 14930 8045 15760 8145 4 S4A
port 1 nsew
rlabel metal2 s 10295 7915 15760 8015 4 S1B
port 2 nsew
rlabel metal2 s 11330 7785 15760 7885 4 S1A
port 3 nsew
rlabel metal2 s 13695 7655 15760 7755 4 S3B
port 4 nsew
rlabel metal2 s 14730 7525 15760 7625 4 S3A
port 5 nsew
rlabel metal2 s 12190 7395 15760 7495 4 S2A
port 6 nsew
rlabel metal2 s 14530 7265 15760 7365 4 S2B
port 7 nsew
rlabel metal2 s 9185 8175 10425 8275 4 S4B
port 8 nsew
rlabel metal2 s 12860 8175 15760 8275 4 S4B
port 8 nsew
rlabel metal2 s 16020 3425 16085 12110 4 BIAS
port 9 nsew
rlabel metal2 s 15925 3760 15990 11765 4 VDD
port 10 nsew
rlabel metal2 s 15825 4175 15890 11400 4 GND
port 11 nsew
rlabel locali s 12290 8660 12670 8695 4 SUB
port 12 nsew
<< end >>
