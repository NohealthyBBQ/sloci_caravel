magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect -5320 3700 -2040 3760
rect -5320 3597 -5220 3700
rect -5320 3563 -5287 3597
rect -5253 3563 -5220 3597
rect -5320 3525 -5220 3563
rect -5320 3491 -5287 3525
rect -5253 3491 -5220 3525
rect -5320 3453 -5220 3491
rect -5320 3419 -5287 3453
rect -5253 3419 -5220 3453
rect -5320 3381 -5220 3419
rect -5320 3347 -5287 3381
rect -5253 3347 -5220 3381
rect -5320 3309 -5220 3347
rect -5320 3275 -5287 3309
rect -5253 3275 -5220 3309
rect -5320 3237 -5220 3275
rect -5320 3203 -5287 3237
rect -5253 3203 -5220 3237
rect -5320 2497 -5220 3203
rect -5320 2463 -5287 2497
rect -5253 2463 -5220 2497
rect -5320 2425 -5220 2463
rect -5320 2391 -5287 2425
rect -5253 2391 -5220 2425
rect -5320 2353 -5220 2391
rect -5320 2319 -5287 2353
rect -5253 2319 -5220 2353
rect -5320 2281 -5220 2319
rect -5320 2247 -5287 2281
rect -5253 2247 -5220 2281
rect -5320 2209 -5220 2247
rect -5320 2175 -5287 2209
rect -5253 2175 -5220 2209
rect -5320 2137 -5220 2175
rect -5320 2103 -5287 2137
rect -5253 2103 -5220 2137
rect -5320 1377 -5220 2103
rect -5320 1343 -5287 1377
rect -5253 1343 -5220 1377
rect -5320 1305 -5220 1343
rect -5320 1271 -5287 1305
rect -5253 1271 -5220 1305
rect -5320 1233 -5220 1271
rect -5320 1199 -5287 1233
rect -5253 1199 -5220 1233
rect -5320 1161 -5220 1199
rect -5320 1127 -5287 1161
rect -5253 1127 -5220 1161
rect -5320 1089 -5220 1127
rect -5320 1055 -5287 1089
rect -5253 1055 -5220 1089
rect -5320 1017 -5220 1055
rect -5320 983 -5287 1017
rect -5253 983 -5220 1017
rect -5320 820 -5220 983
rect -4080 900 -4000 3700
rect -4080 820 -2040 900
rect 4820 837 5140 860
rect 4820 803 4855 837
rect 4889 803 4927 837
rect 4961 803 4999 837
rect 5033 803 5071 837
rect 5105 803 5140 837
rect 4820 780 5140 803
<< viali >>
rect -5287 3563 -5253 3597
rect -5287 3491 -5253 3525
rect -5287 3419 -5253 3453
rect -5287 3347 -5253 3381
rect -5287 3275 -5253 3309
rect -5287 3203 -5253 3237
rect -5287 2463 -5253 2497
rect -5287 2391 -5253 2425
rect -5287 2319 -5253 2353
rect -5287 2247 -5253 2281
rect -5287 2175 -5253 2209
rect -5287 2103 -5253 2137
rect -5287 1343 -5253 1377
rect -5287 1271 -5253 1305
rect -5287 1199 -5253 1233
rect -5287 1127 -5253 1161
rect -5287 1055 -5253 1089
rect -5287 983 -5253 1017
rect 4855 803 4889 837
rect 4927 803 4961 837
rect 4999 803 5033 837
rect 5071 803 5105 837
<< metal1 >>
rect -5170 5676 -4750 5680
rect -5170 5624 -5146 5676
rect -5094 5624 -5082 5676
rect -5030 5624 -5018 5676
rect -4966 5624 -4954 5676
rect -4902 5624 -4890 5676
rect -4838 5624 -4826 5676
rect -4774 5624 -4750 5676
rect -5170 5620 -4750 5624
rect -3730 5676 -3310 5680
rect -3730 5624 -3706 5676
rect -3654 5624 -3642 5676
rect -3590 5624 -3578 5676
rect -3526 5624 -3514 5676
rect -3462 5624 -3450 5676
rect -3398 5624 -3386 5676
rect -3334 5624 -3310 5676
rect -3730 5620 -3310 5624
rect -2690 5676 -2270 5680
rect -2690 5624 -2666 5676
rect -2614 5624 -2602 5676
rect -2550 5624 -2538 5676
rect -2486 5624 -2474 5676
rect -2422 5624 -2410 5676
rect -2358 5624 -2346 5676
rect -2294 5624 -2270 5676
rect -2690 5620 -2270 5624
rect -1230 5676 -810 5680
rect -1230 5624 -1206 5676
rect -1154 5624 -1142 5676
rect -1090 5624 -1078 5676
rect -1026 5624 -1014 5676
rect -962 5624 -950 5676
rect -898 5624 -886 5676
rect -834 5624 -810 5676
rect -1230 5620 -810 5624
rect -5170 4096 -4750 4100
rect -5170 4044 -5146 4096
rect -5094 4044 -5082 4096
rect -5030 4044 -5018 4096
rect -4966 4044 -4954 4096
rect -4902 4044 -4890 4096
rect -4838 4044 -4826 4096
rect -4774 4044 -4750 4096
rect -3730 4044 -3720 4100
rect -3320 4044 -3310 4100
rect -2272 4044 -2270 4100
rect -1230 4096 -810 4100
rect -1230 4044 -1206 4096
rect -1154 4044 -1142 4096
rect -1090 4044 -1078 4096
rect -1026 4044 -1014 4096
rect -962 4044 -950 4096
rect -898 4044 -886 4096
rect -834 4044 -810 4096
rect -5170 4040 -4750 4044
rect -1230 4040 -810 4044
rect -5306 3600 -5234 3612
rect -5310 3597 -5230 3600
rect -5310 3586 -5287 3597
rect -5253 3586 -5230 3597
rect -5310 3534 -5296 3586
rect -5244 3534 -5230 3586
rect -5310 3525 -5230 3534
rect -5310 3522 -5287 3525
rect -5253 3522 -5230 3525
rect -5310 3470 -5296 3522
rect -5244 3470 -5230 3522
rect -5310 3458 -5230 3470
rect -5310 3406 -5296 3458
rect -5244 3406 -5230 3458
rect -5310 3394 -5230 3406
rect -5310 3342 -5296 3394
rect -5244 3342 -5230 3394
rect -5310 3330 -5230 3342
rect -5310 3278 -5296 3330
rect -5244 3278 -5230 3330
rect -5310 3275 -5287 3278
rect -5253 3275 -5230 3278
rect -5310 3266 -5230 3275
rect -5310 3214 -5296 3266
rect -5244 3214 -5230 3266
rect -5310 3203 -5287 3214
rect -5253 3203 -5230 3214
rect -5310 3200 -5230 3203
rect -4100 3226 -3980 3720
rect -5306 3188 -5234 3200
rect -4100 3174 -4056 3226
rect -4004 3174 -3980 3226
rect -4100 3162 -3980 3174
rect -4100 3110 -4056 3162
rect -4004 3110 -3980 3162
rect -4100 3098 -3980 3110
rect -4100 3046 -4056 3098
rect -4004 3046 -3980 3098
rect -4100 3034 -3980 3046
rect -4100 2982 -4056 3034
rect -4004 2982 -3980 3034
rect -4100 2970 -3980 2982
rect -4100 2918 -4056 2970
rect -4004 2918 -3980 2970
rect -4100 2906 -3980 2918
rect -4100 2854 -4056 2906
rect -4004 2854 -3980 2906
rect -5306 2500 -5234 2512
rect -5310 2497 -5230 2500
rect -5310 2486 -5287 2497
rect -5253 2486 -5230 2497
rect -5310 2434 -5296 2486
rect -5244 2434 -5230 2486
rect -5310 2425 -5230 2434
rect -5310 2422 -5287 2425
rect -5253 2422 -5230 2425
rect -5310 2370 -5296 2422
rect -5244 2370 -5230 2422
rect -5310 2358 -5230 2370
rect -5310 2306 -5296 2358
rect -5244 2306 -5230 2358
rect -5310 2294 -5230 2306
rect -5310 2242 -5296 2294
rect -5244 2242 -5230 2294
rect -5310 2230 -5230 2242
rect -5310 2178 -5296 2230
rect -5244 2178 -5230 2230
rect -5310 2175 -5287 2178
rect -5253 2175 -5230 2178
rect -5310 2166 -5230 2175
rect -5310 2114 -5296 2166
rect -5244 2114 -5230 2166
rect -5310 2103 -5287 2114
rect -5253 2103 -5230 2114
rect -5310 2100 -5230 2103
rect -4100 2106 -3980 2854
rect 510 2656 590 2660
rect 510 2604 524 2656
rect 576 2604 590 2656
rect 510 2600 590 2604
rect -5306 2088 -5234 2100
rect -4100 2054 -4056 2106
rect -4004 2054 -3980 2106
rect -4100 2042 -3980 2054
rect -4100 1990 -4056 2042
rect -4004 1990 -3980 2042
rect -4100 1978 -3980 1990
rect -4100 1926 -4056 1978
rect -4004 1926 -3980 1978
rect -4100 1914 -3980 1926
rect -4100 1862 -4056 1914
rect -4004 1862 -3980 1914
rect -4100 1850 -3980 1862
rect -4100 1798 -4056 1850
rect -4004 1798 -3980 1850
rect -4100 1786 -3980 1798
rect -4100 1734 -4056 1786
rect -4004 1734 -3980 1786
rect -5306 1380 -5234 1392
rect -5310 1377 -5230 1380
rect -5310 1366 -5287 1377
rect -5253 1366 -5230 1377
rect -5310 1314 -5296 1366
rect -5244 1314 -5230 1366
rect -5310 1305 -5230 1314
rect -5310 1302 -5287 1305
rect -5253 1302 -5230 1305
rect -5310 1250 -5296 1302
rect -5244 1250 -5230 1302
rect -5310 1238 -5230 1250
rect -5310 1186 -5296 1238
rect -5244 1186 -5230 1238
rect -5310 1174 -5230 1186
rect -5310 1122 -5296 1174
rect -5244 1122 -5230 1174
rect -5310 1110 -5230 1122
rect -5310 1058 -5296 1110
rect -5244 1058 -5230 1110
rect -5310 1055 -5287 1058
rect -5253 1055 -5230 1058
rect -5310 1046 -5230 1055
rect -5310 994 -5296 1046
rect -5244 994 -5230 1046
rect -5310 983 -5287 994
rect -5253 983 -5230 994
rect -5310 980 -5230 983
rect -5306 968 -5234 980
rect -4685 770 -4625 966
rect -4100 880 -3980 1734
rect 6290 1372 6510 1400
rect 6290 1128 6310 1372
rect 6490 1128 6510 1372
rect 6290 1100 6510 1128
rect 3346 1005 3441 1031
rect 3346 966 3367 1005
rect 3338 953 3367 966
rect 3419 963 3441 1005
rect 3419 953 3459 963
rect -3470 936 -2750 940
rect -3470 884 -3456 936
rect -3404 884 -3392 936
rect -3340 884 -3328 936
rect -3276 884 -3264 936
rect -3212 884 -3200 936
rect -3148 884 -3136 936
rect -3084 884 -3072 936
rect -3020 884 -3008 936
rect -2956 884 -2944 936
rect -2892 884 -2880 936
rect -2828 884 -2816 936
rect -2764 884 -2750 936
rect 3338 907 3459 953
rect -3470 880 -2750 884
rect 4808 846 5152 866
rect 4808 794 4826 846
rect 4878 837 4890 846
rect 4942 837 4954 846
rect 5006 837 5018 846
rect 5070 837 5082 846
rect 4889 803 4890 837
rect 5070 803 5071 837
rect 4878 794 4890 803
rect 4942 794 4954 803
rect 5006 794 5018 803
rect 5070 794 5082 803
rect 5134 794 5152 846
rect 4808 774 5152 794
rect -4685 710 -750 770
rect -4685 701 -4625 710
rect -1324 594 -1276 710
<< via1 >>
rect -5146 5624 -5094 5676
rect -5082 5624 -5030 5676
rect -5018 5624 -4966 5676
rect -4954 5624 -4902 5676
rect -4890 5624 -4838 5676
rect -4826 5624 -4774 5676
rect -3706 5624 -3654 5676
rect -3642 5624 -3590 5676
rect -3578 5624 -3526 5676
rect -3514 5624 -3462 5676
rect -3450 5624 -3398 5676
rect -3386 5624 -3334 5676
rect -2666 5624 -2614 5676
rect -2602 5624 -2550 5676
rect -2538 5624 -2486 5676
rect -2474 5624 -2422 5676
rect -2410 5624 -2358 5676
rect -2346 5624 -2294 5676
rect -1206 5624 -1154 5676
rect -1142 5624 -1090 5676
rect -1078 5624 -1026 5676
rect -1014 5624 -962 5676
rect -950 5624 -898 5676
rect -886 5624 -834 5676
rect -5146 4044 -5094 4096
rect -5082 4044 -5030 4096
rect -5018 4044 -4966 4096
rect -4954 4044 -4902 4096
rect -4890 4044 -4838 4096
rect -4826 4044 -4774 4096
rect -1206 4044 -1154 4096
rect -1142 4044 -1090 4096
rect -1078 4044 -1026 4096
rect -1014 4044 -962 4096
rect -950 4044 -898 4096
rect -886 4044 -834 4096
rect -5296 3563 -5287 3586
rect -5287 3563 -5253 3586
rect -5253 3563 -5244 3586
rect -5296 3534 -5244 3563
rect -5296 3491 -5287 3522
rect -5287 3491 -5253 3522
rect -5253 3491 -5244 3522
rect -5296 3470 -5244 3491
rect -5296 3453 -5244 3458
rect -5296 3419 -5287 3453
rect -5287 3419 -5253 3453
rect -5253 3419 -5244 3453
rect -5296 3406 -5244 3419
rect -5296 3381 -5244 3394
rect -5296 3347 -5287 3381
rect -5287 3347 -5253 3381
rect -5253 3347 -5244 3381
rect -5296 3342 -5244 3347
rect -5296 3309 -5244 3330
rect -5296 3278 -5287 3309
rect -5287 3278 -5253 3309
rect -5253 3278 -5244 3309
rect -5296 3237 -5244 3266
rect -5296 3214 -5287 3237
rect -5287 3214 -5253 3237
rect -5253 3214 -5244 3237
rect -4056 3174 -4004 3226
rect -4056 3110 -4004 3162
rect -4056 3046 -4004 3098
rect -4056 2982 -4004 3034
rect -4056 2918 -4004 2970
rect -4056 2854 -4004 2906
rect -5296 2463 -5287 2486
rect -5287 2463 -5253 2486
rect -5253 2463 -5244 2486
rect -5296 2434 -5244 2463
rect -5296 2391 -5287 2422
rect -5287 2391 -5253 2422
rect -5253 2391 -5244 2422
rect -5296 2370 -5244 2391
rect -5296 2353 -5244 2358
rect -5296 2319 -5287 2353
rect -5287 2319 -5253 2353
rect -5253 2319 -5244 2353
rect -5296 2306 -5244 2319
rect -5296 2281 -5244 2294
rect -5296 2247 -5287 2281
rect -5287 2247 -5253 2281
rect -5253 2247 -5244 2281
rect -5296 2242 -5244 2247
rect -5296 2209 -5244 2230
rect -5296 2178 -5287 2209
rect -5287 2178 -5253 2209
rect -5253 2178 -5244 2209
rect -5296 2137 -5244 2166
rect -5296 2114 -5287 2137
rect -5287 2114 -5253 2137
rect -5253 2114 -5244 2137
rect 524 2604 576 2656
rect -4056 2054 -4004 2106
rect -4056 1990 -4004 2042
rect -4056 1926 -4004 1978
rect -4056 1862 -4004 1914
rect -4056 1798 -4004 1850
rect -4056 1734 -4004 1786
rect -5296 1343 -5287 1366
rect -5287 1343 -5253 1366
rect -5253 1343 -5244 1366
rect -5296 1314 -5244 1343
rect -5296 1271 -5287 1302
rect -5287 1271 -5253 1302
rect -5253 1271 -5244 1302
rect -5296 1250 -5244 1271
rect -5296 1233 -5244 1238
rect -5296 1199 -5287 1233
rect -5287 1199 -5253 1233
rect -5253 1199 -5244 1233
rect -5296 1186 -5244 1199
rect -5296 1161 -5244 1174
rect -5296 1127 -5287 1161
rect -5287 1127 -5253 1161
rect -5253 1127 -5244 1161
rect -5296 1122 -5244 1127
rect -5296 1089 -5244 1110
rect -5296 1058 -5287 1089
rect -5287 1058 -5253 1089
rect -5253 1058 -5244 1089
rect -5296 1017 -5244 1046
rect -5296 994 -5287 1017
rect -5287 994 -5253 1017
rect -5253 994 -5244 1017
rect 6310 1128 6490 1372
rect 3367 953 3419 1005
rect -3456 884 -3404 936
rect -3392 884 -3340 936
rect -3328 884 -3276 936
rect -3264 884 -3212 936
rect -3200 884 -3148 936
rect -3136 884 -3084 936
rect -3072 884 -3020 936
rect -3008 884 -2956 936
rect -2944 884 -2892 936
rect -2880 884 -2828 936
rect -2816 884 -2764 936
rect 4826 837 4878 846
rect 4890 837 4942 846
rect 4954 837 5006 846
rect 5018 837 5070 846
rect 5082 837 5134 846
rect 4826 803 4855 837
rect 4855 803 4878 837
rect 4890 803 4927 837
rect 4927 803 4942 837
rect 4954 803 4961 837
rect 4961 803 4999 837
rect 4999 803 5006 837
rect 5018 803 5033 837
rect 5033 803 5070 837
rect 5082 803 5105 837
rect 5105 803 5134 837
rect 4826 794 4878 803
rect 4890 794 4942 803
rect 4954 794 5006 803
rect 5018 794 5070 803
rect 5082 794 5134 803
<< metal2 >>
rect -5160 5678 -4760 5690
rect -5160 5622 -5148 5678
rect -5092 5676 -5068 5678
rect -5012 5676 -4988 5678
rect -4932 5676 -4908 5678
rect -4852 5676 -4828 5678
rect -5092 5624 -5082 5676
rect -4838 5624 -4828 5676
rect -5092 5622 -5068 5624
rect -5012 5622 -4988 5624
rect -4932 5622 -4908 5624
rect -4852 5622 -4828 5624
rect -4772 5622 -4760 5678
rect -5160 5610 -4760 5622
rect -3720 5678 -3320 5690
rect -3720 5622 -3708 5678
rect -3652 5676 -3628 5678
rect -3572 5676 -3548 5678
rect -3492 5676 -3468 5678
rect -3412 5676 -3388 5678
rect -3652 5624 -3642 5676
rect -3398 5624 -3388 5676
rect -3652 5622 -3628 5624
rect -3572 5622 -3548 5624
rect -3492 5622 -3468 5624
rect -3412 5622 -3388 5624
rect -3332 5622 -3320 5678
rect -3720 5610 -3320 5622
rect -2680 5678 -2280 5690
rect -2680 5622 -2668 5678
rect -2612 5676 -2588 5678
rect -2532 5676 -2508 5678
rect -2452 5676 -2428 5678
rect -2372 5676 -2348 5678
rect -2612 5624 -2602 5676
rect -2358 5624 -2348 5676
rect -2612 5622 -2588 5624
rect -2532 5622 -2508 5624
rect -2452 5622 -2428 5624
rect -2372 5622 -2348 5624
rect -2292 5622 -2280 5678
rect -2680 5610 -2280 5622
rect -1220 5678 -820 5690
rect -1220 5622 -1208 5678
rect -1152 5676 -1128 5678
rect -1072 5676 -1048 5678
rect -992 5676 -968 5678
rect -912 5676 -888 5678
rect -1152 5624 -1142 5676
rect -898 5624 -888 5676
rect -1152 5622 -1128 5624
rect -1072 5622 -1048 5624
rect -992 5622 -968 5624
rect -912 5622 -888 5624
rect -832 5622 -820 5678
rect -1220 5610 -820 5622
rect -5160 4098 -4760 4110
rect -5160 4042 -5148 4098
rect -5092 4096 -5068 4098
rect -5012 4096 -4988 4098
rect -4932 4096 -4908 4098
rect -4852 4096 -4828 4098
rect -5092 4044 -5082 4096
rect -4838 4044 -4828 4096
rect -5092 4042 -5068 4044
rect -5012 4042 -4988 4044
rect -4932 4042 -4908 4044
rect -4852 4042 -4828 4044
rect -4772 4042 -4760 4098
rect -5160 4030 -4760 4042
rect -1220 4098 -820 4110
rect -1220 4042 -1208 4098
rect -1152 4096 -1128 4098
rect -1072 4096 -1048 4098
rect -992 4096 -968 4098
rect -912 4096 -888 4098
rect -1152 4044 -1142 4096
rect -898 4044 -888 4096
rect -1152 4042 -1128 4044
rect -1072 4042 -1048 4044
rect -992 4042 -968 4044
rect -912 4042 -888 4044
rect -832 4042 -820 4098
rect -1220 4030 -820 4042
rect 300 3670 650 3800
rect -5300 3588 -5240 3610
rect -5300 3532 -5298 3588
rect -5242 3532 -5240 3588
rect -5300 3522 -5240 3532
rect -5300 3508 -5296 3522
rect -5244 3508 -5240 3522
rect -5300 3452 -5298 3508
rect -5242 3452 -5240 3508
rect -5300 3428 -5296 3452
rect -5244 3428 -5240 3452
rect -5300 3372 -5298 3428
rect -5242 3372 -5240 3428
rect -5300 3348 -5296 3372
rect -5244 3348 -5240 3372
rect -5300 3292 -5298 3348
rect -5242 3292 -5240 3348
rect -5300 3278 -5296 3292
rect -5244 3278 -5240 3292
rect -5300 3268 -5240 3278
rect -5300 3212 -5298 3268
rect -5242 3212 -5240 3268
rect -5300 3190 -5240 3212
rect -4060 3228 -4000 3250
rect -4060 3172 -4058 3228
rect -4002 3172 -4000 3228
rect -4060 3162 -4000 3172
rect -4060 3148 -4056 3162
rect -4004 3148 -4000 3162
rect -4060 3092 -4058 3148
rect -4002 3092 -4000 3148
rect -4060 3068 -4056 3092
rect -4004 3068 -4000 3092
rect -4060 3012 -4058 3068
rect -4002 3012 -4000 3068
rect -4060 2988 -4056 3012
rect -4004 2988 -4000 3012
rect -4060 2932 -4058 2988
rect -4002 2932 -4000 2988
rect -4060 2918 -4056 2932
rect -4004 2918 -4000 2932
rect -4060 2908 -4000 2918
rect 280 2913 736 3045
rect -4060 2852 -4058 2908
rect -4002 2852 -4000 2908
rect -4060 2830 -4000 2852
rect -3780 2658 -3710 2670
rect -3780 2602 -3773 2658
rect -3717 2602 -3710 2658
rect -3780 2590 -3710 2602
rect -2480 2658 590 2670
rect -2480 2602 -1733 2658
rect -1677 2656 590 2658
rect -1677 2604 524 2656
rect 576 2604 590 2656
rect -1677 2602 590 2604
rect -2480 2590 590 2602
rect -5300 2488 -5240 2510
rect -5300 2432 -5298 2488
rect -5242 2432 -5240 2488
rect -5300 2422 -5240 2432
rect -5300 2408 -5296 2422
rect -5244 2408 -5240 2422
rect -5300 2352 -5298 2408
rect -5242 2352 -5240 2408
rect -2752 2352 -2652 2432
rect -5300 2328 -5296 2352
rect -5244 2328 -5240 2352
rect -5300 2272 -5298 2328
rect -5242 2272 -5240 2328
rect -5300 2248 -5296 2272
rect -5244 2248 -5240 2272
rect -4080 2328 -4000 2340
rect -4080 2272 -4068 2328
rect -4012 2272 -4000 2328
rect -4080 2260 -4000 2272
rect -5300 2192 -5298 2248
rect -5242 2192 -5240 2248
rect -5300 2178 -5296 2192
rect -5244 2178 -5240 2192
rect -5300 2168 -5240 2178
rect -2752 2172 -2652 2252
rect -5300 2112 -5298 2168
rect -5242 2112 -5240 2168
rect 301 2157 647 2289
rect -5300 2090 -5240 2112
rect -4060 2108 -4000 2130
rect -4060 2052 -4058 2108
rect -4002 2052 -4000 2108
rect -4060 2042 -4000 2052
rect -4060 2028 -4056 2042
rect -4004 2028 -4000 2042
rect -4060 1972 -4058 2028
rect -4002 1972 -4000 2028
rect -4060 1948 -4056 1972
rect -4004 1948 -4000 1972
rect -4060 1892 -4058 1948
rect -4002 1892 -4000 1948
rect -4060 1868 -4056 1892
rect -4004 1868 -4000 1892
rect -4060 1812 -4058 1868
rect -4002 1812 -4000 1868
rect -4060 1798 -4056 1812
rect -4004 1798 -4000 1812
rect -4060 1788 -4000 1798
rect -4060 1732 -4058 1788
rect -4002 1732 -4000 1788
rect -4060 1710 -4000 1732
rect 305 1401 651 1533
rect 6300 1398 6500 1410
rect -5300 1368 -5240 1390
rect -5300 1312 -5298 1368
rect -5242 1312 -5240 1368
rect -5300 1302 -5240 1312
rect -5300 1288 -5296 1302
rect -5244 1288 -5240 1302
rect -5300 1232 -5298 1288
rect -5242 1232 -5240 1288
rect -5300 1208 -5296 1232
rect -5244 1208 -5240 1232
rect -5300 1152 -5298 1208
rect -5242 1152 -5240 1208
rect -5300 1128 -5296 1152
rect -5244 1128 -5240 1152
rect -5300 1072 -5298 1128
rect -5242 1072 -5240 1128
rect 6300 1372 6332 1398
rect 6468 1372 6500 1398
rect 6300 1128 6310 1372
rect 6490 1128 6500 1372
rect 6300 1102 6332 1128
rect 6468 1102 6500 1128
rect 6300 1090 6500 1102
rect -5300 1058 -5296 1072
rect -5244 1058 -5240 1072
rect -5300 1048 -5240 1058
rect -5300 992 -5298 1048
rect -5242 992 -5240 1048
rect -5300 970 -5240 992
rect 3009 1005 3459 1047
rect 3009 953 3367 1005
rect 3419 953 3459 1005
rect -3460 936 -2760 950
rect -3460 884 -3456 936
rect -3404 884 -3392 936
rect -3340 884 -3328 936
rect -3276 884 -3264 936
rect -3212 884 -3200 936
rect -3148 884 -3136 936
rect -3084 884 -3072 936
rect -3020 884 -3008 936
rect -2956 884 -2944 936
rect -2892 884 -2880 936
rect -2828 884 -2816 936
rect -2764 884 -2760 936
rect 3009 907 3459 953
rect -3460 798 -2760 884
rect -3460 742 -3458 798
rect -3402 742 -3378 798
rect -3322 742 -3298 798
rect -3242 742 -3218 798
rect -3162 742 -3138 798
rect -3082 742 -3058 798
rect -3002 742 -2978 798
rect -2922 742 -2898 798
rect -2842 742 -2818 798
rect -2762 742 -2760 798
rect 4820 848 5140 870
rect 4820 846 4832 848
rect 4888 846 4912 848
rect 4968 846 4992 848
rect 5048 846 5072 848
rect 5128 846 5140 848
rect 4820 794 4826 846
rect 4888 794 4890 846
rect 5070 794 5072 846
rect 5134 794 5140 846
rect 4820 792 4832 794
rect 4888 792 4912 794
rect 4968 792 4992 794
rect 5048 792 5072 794
rect 5128 792 5140 794
rect 4820 770 5140 792
rect -3460 730 -2760 742
<< via2 >>
rect -5148 5676 -5092 5678
rect -5068 5676 -5012 5678
rect -4988 5676 -4932 5678
rect -4908 5676 -4852 5678
rect -4828 5676 -4772 5678
rect -5148 5624 -5146 5676
rect -5146 5624 -5094 5676
rect -5094 5624 -5092 5676
rect -5068 5624 -5030 5676
rect -5030 5624 -5018 5676
rect -5018 5624 -5012 5676
rect -4988 5624 -4966 5676
rect -4966 5624 -4954 5676
rect -4954 5624 -4932 5676
rect -4908 5624 -4902 5676
rect -4902 5624 -4890 5676
rect -4890 5624 -4852 5676
rect -4828 5624 -4826 5676
rect -4826 5624 -4774 5676
rect -4774 5624 -4772 5676
rect -5148 5622 -5092 5624
rect -5068 5622 -5012 5624
rect -4988 5622 -4932 5624
rect -4908 5622 -4852 5624
rect -4828 5622 -4772 5624
rect -3708 5676 -3652 5678
rect -3628 5676 -3572 5678
rect -3548 5676 -3492 5678
rect -3468 5676 -3412 5678
rect -3388 5676 -3332 5678
rect -3708 5624 -3706 5676
rect -3706 5624 -3654 5676
rect -3654 5624 -3652 5676
rect -3628 5624 -3590 5676
rect -3590 5624 -3578 5676
rect -3578 5624 -3572 5676
rect -3548 5624 -3526 5676
rect -3526 5624 -3514 5676
rect -3514 5624 -3492 5676
rect -3468 5624 -3462 5676
rect -3462 5624 -3450 5676
rect -3450 5624 -3412 5676
rect -3388 5624 -3386 5676
rect -3386 5624 -3334 5676
rect -3334 5624 -3332 5676
rect -3708 5622 -3652 5624
rect -3628 5622 -3572 5624
rect -3548 5622 -3492 5624
rect -3468 5622 -3412 5624
rect -3388 5622 -3332 5624
rect -2668 5676 -2612 5678
rect -2588 5676 -2532 5678
rect -2508 5676 -2452 5678
rect -2428 5676 -2372 5678
rect -2348 5676 -2292 5678
rect -2668 5624 -2666 5676
rect -2666 5624 -2614 5676
rect -2614 5624 -2612 5676
rect -2588 5624 -2550 5676
rect -2550 5624 -2538 5676
rect -2538 5624 -2532 5676
rect -2508 5624 -2486 5676
rect -2486 5624 -2474 5676
rect -2474 5624 -2452 5676
rect -2428 5624 -2422 5676
rect -2422 5624 -2410 5676
rect -2410 5624 -2372 5676
rect -2348 5624 -2346 5676
rect -2346 5624 -2294 5676
rect -2294 5624 -2292 5676
rect -2668 5622 -2612 5624
rect -2588 5622 -2532 5624
rect -2508 5622 -2452 5624
rect -2428 5622 -2372 5624
rect -2348 5622 -2292 5624
rect -1208 5676 -1152 5678
rect -1128 5676 -1072 5678
rect -1048 5676 -992 5678
rect -968 5676 -912 5678
rect -888 5676 -832 5678
rect -1208 5624 -1206 5676
rect -1206 5624 -1154 5676
rect -1154 5624 -1152 5676
rect -1128 5624 -1090 5676
rect -1090 5624 -1078 5676
rect -1078 5624 -1072 5676
rect -1048 5624 -1026 5676
rect -1026 5624 -1014 5676
rect -1014 5624 -992 5676
rect -968 5624 -962 5676
rect -962 5624 -950 5676
rect -950 5624 -912 5676
rect -888 5624 -886 5676
rect -886 5624 -834 5676
rect -834 5624 -832 5676
rect -1208 5622 -1152 5624
rect -1128 5622 -1072 5624
rect -1048 5622 -992 5624
rect -968 5622 -912 5624
rect -888 5622 -832 5624
rect -5148 4096 -5092 4098
rect -5068 4096 -5012 4098
rect -4988 4096 -4932 4098
rect -4908 4096 -4852 4098
rect -4828 4096 -4772 4098
rect -5148 4044 -5146 4096
rect -5146 4044 -5094 4096
rect -5094 4044 -5092 4096
rect -5068 4044 -5030 4096
rect -5030 4044 -5018 4096
rect -5018 4044 -5012 4096
rect -4988 4044 -4966 4096
rect -4966 4044 -4954 4096
rect -4954 4044 -4932 4096
rect -4908 4044 -4902 4096
rect -4902 4044 -4890 4096
rect -4890 4044 -4852 4096
rect -4828 4044 -4826 4096
rect -4826 4044 -4774 4096
rect -4774 4044 -4772 4096
rect -5148 4042 -5092 4044
rect -5068 4042 -5012 4044
rect -4988 4042 -4932 4044
rect -4908 4042 -4852 4044
rect -4828 4042 -4772 4044
rect -1208 4096 -1152 4098
rect -1128 4096 -1072 4098
rect -1048 4096 -992 4098
rect -968 4096 -912 4098
rect -888 4096 -832 4098
rect -1208 4044 -1206 4096
rect -1206 4044 -1154 4096
rect -1154 4044 -1152 4096
rect -1128 4044 -1090 4096
rect -1090 4044 -1078 4096
rect -1078 4044 -1072 4096
rect -1048 4044 -1026 4096
rect -1026 4044 -1014 4096
rect -1014 4044 -992 4096
rect -968 4044 -962 4096
rect -962 4044 -950 4096
rect -950 4044 -912 4096
rect -888 4044 -886 4096
rect -886 4044 -834 4096
rect -834 4044 -832 4096
rect -1208 4042 -1152 4044
rect -1128 4042 -1072 4044
rect -1048 4042 -992 4044
rect -968 4042 -912 4044
rect -888 4042 -832 4044
rect -5298 3586 -5242 3588
rect -5298 3534 -5296 3586
rect -5296 3534 -5244 3586
rect -5244 3534 -5242 3586
rect -5298 3532 -5242 3534
rect -5298 3470 -5296 3508
rect -5296 3470 -5244 3508
rect -5244 3470 -5242 3508
rect -5298 3458 -5242 3470
rect -5298 3452 -5296 3458
rect -5296 3452 -5244 3458
rect -5244 3452 -5242 3458
rect -5298 3406 -5296 3428
rect -5296 3406 -5244 3428
rect -5244 3406 -5242 3428
rect -5298 3394 -5242 3406
rect -5298 3372 -5296 3394
rect -5296 3372 -5244 3394
rect -5244 3372 -5242 3394
rect -5298 3342 -5296 3348
rect -5296 3342 -5244 3348
rect -5244 3342 -5242 3348
rect -5298 3330 -5242 3342
rect -5298 3292 -5296 3330
rect -5296 3292 -5244 3330
rect -5244 3292 -5242 3330
rect -5298 3266 -5242 3268
rect -5298 3214 -5296 3266
rect -5296 3214 -5244 3266
rect -5244 3214 -5242 3266
rect -5298 3212 -5242 3214
rect -4058 3226 -4002 3228
rect -4058 3174 -4056 3226
rect -4056 3174 -4004 3226
rect -4004 3174 -4002 3226
rect -4058 3172 -4002 3174
rect -4058 3110 -4056 3148
rect -4056 3110 -4004 3148
rect -4004 3110 -4002 3148
rect -4058 3098 -4002 3110
rect -4058 3092 -4056 3098
rect -4056 3092 -4004 3098
rect -4004 3092 -4002 3098
rect -4058 3046 -4056 3068
rect -4056 3046 -4004 3068
rect -4004 3046 -4002 3068
rect -4058 3034 -4002 3046
rect -4058 3012 -4056 3034
rect -4056 3012 -4004 3034
rect -4004 3012 -4002 3034
rect -4058 2982 -4056 2988
rect -4056 2982 -4004 2988
rect -4004 2982 -4002 2988
rect -4058 2970 -4002 2982
rect -4058 2932 -4056 2970
rect -4056 2932 -4004 2970
rect -4004 2932 -4002 2970
rect -4058 2906 -4002 2908
rect -4058 2854 -4056 2906
rect -4056 2854 -4004 2906
rect -4004 2854 -4002 2906
rect -4058 2852 -4002 2854
rect -3773 2602 -3717 2658
rect -1733 2602 -1677 2658
rect -5298 2486 -5242 2488
rect -5298 2434 -5296 2486
rect -5296 2434 -5244 2486
rect -5244 2434 -5242 2486
rect -5298 2432 -5242 2434
rect -5298 2370 -5296 2408
rect -5296 2370 -5244 2408
rect -5244 2370 -5242 2408
rect -5298 2358 -5242 2370
rect -5298 2352 -5296 2358
rect -5296 2352 -5244 2358
rect -5244 2352 -5242 2358
rect -5298 2306 -5296 2328
rect -5296 2306 -5244 2328
rect -5244 2306 -5242 2328
rect -5298 2294 -5242 2306
rect -5298 2272 -5296 2294
rect -5296 2272 -5244 2294
rect -5244 2272 -5242 2294
rect -4068 2272 -4012 2328
rect -5298 2242 -5296 2248
rect -5296 2242 -5244 2248
rect -5244 2242 -5242 2248
rect -5298 2230 -5242 2242
rect -5298 2192 -5296 2230
rect -5296 2192 -5244 2230
rect -5244 2192 -5242 2230
rect -5298 2166 -5242 2168
rect -5298 2114 -5296 2166
rect -5296 2114 -5244 2166
rect -5244 2114 -5242 2166
rect -5298 2112 -5242 2114
rect -4058 2106 -4002 2108
rect -4058 2054 -4056 2106
rect -4056 2054 -4004 2106
rect -4004 2054 -4002 2106
rect -4058 2052 -4002 2054
rect -4058 1990 -4056 2028
rect -4056 1990 -4004 2028
rect -4004 1990 -4002 2028
rect -4058 1978 -4002 1990
rect -4058 1972 -4056 1978
rect -4056 1972 -4004 1978
rect -4004 1972 -4002 1978
rect -4058 1926 -4056 1948
rect -4056 1926 -4004 1948
rect -4004 1926 -4002 1948
rect -4058 1914 -4002 1926
rect -4058 1892 -4056 1914
rect -4056 1892 -4004 1914
rect -4004 1892 -4002 1914
rect -4058 1862 -4056 1868
rect -4056 1862 -4004 1868
rect -4004 1862 -4002 1868
rect -4058 1850 -4002 1862
rect -4058 1812 -4056 1850
rect -4056 1812 -4004 1850
rect -4004 1812 -4002 1850
rect -4058 1786 -4002 1788
rect -4058 1734 -4056 1786
rect -4056 1734 -4004 1786
rect -4004 1734 -4002 1786
rect -4058 1732 -4002 1734
rect -5298 1366 -5242 1368
rect -5298 1314 -5296 1366
rect -5296 1314 -5244 1366
rect -5244 1314 -5242 1366
rect -5298 1312 -5242 1314
rect -5298 1250 -5296 1288
rect -5296 1250 -5244 1288
rect -5244 1250 -5242 1288
rect -5298 1238 -5242 1250
rect -5298 1232 -5296 1238
rect -5296 1232 -5244 1238
rect -5244 1232 -5242 1238
rect -5298 1186 -5296 1208
rect -5296 1186 -5244 1208
rect -5244 1186 -5242 1208
rect -5298 1174 -5242 1186
rect -5298 1152 -5296 1174
rect -5296 1152 -5244 1174
rect -5244 1152 -5242 1174
rect -5298 1122 -5296 1128
rect -5296 1122 -5244 1128
rect -5244 1122 -5242 1128
rect -5298 1110 -5242 1122
rect -5298 1072 -5296 1110
rect -5296 1072 -5244 1110
rect -5244 1072 -5242 1110
rect 6332 1372 6468 1398
rect 6332 1128 6468 1372
rect 6332 1102 6468 1128
rect -5298 1046 -5242 1048
rect -5298 994 -5296 1046
rect -5296 994 -5244 1046
rect -5244 994 -5242 1046
rect -5298 992 -5242 994
rect -3458 742 -3402 798
rect -3378 742 -3322 798
rect -3298 742 -3242 798
rect -3218 742 -3162 798
rect -3138 742 -3082 798
rect -3058 742 -3002 798
rect -2978 742 -2922 798
rect -2898 742 -2842 798
rect -2818 742 -2762 798
rect 4832 846 4888 848
rect 4912 846 4968 848
rect 4992 846 5048 848
rect 5072 846 5128 848
rect 4832 794 4878 846
rect 4878 794 4888 846
rect 4912 794 4942 846
rect 4942 794 4954 846
rect 4954 794 4968 846
rect 4992 794 5006 846
rect 5006 794 5018 846
rect 5018 794 5048 846
rect 5072 794 5082 846
rect 5082 794 5128 846
rect 4832 792 4888 794
rect 4912 792 4968 794
rect 4992 792 5048 794
rect 5072 792 5128 794
<< metal3 >>
rect 1810 5772 1950 5780
rect -5170 5702 -4750 5720
rect -5170 5638 -5152 5702
rect -5088 5638 -5072 5702
rect -5008 5638 -4992 5702
rect -4928 5638 -4912 5702
rect -4848 5638 -4832 5702
rect -4768 5638 -4750 5702
rect -5170 5622 -5148 5638
rect -5092 5622 -5068 5638
rect -5012 5622 -4988 5638
rect -4932 5622 -4908 5638
rect -4852 5622 -4828 5638
rect -4772 5622 -4750 5638
rect -5170 5615 -4750 5622
rect -3730 5702 -3310 5720
rect -3730 5638 -3712 5702
rect -3648 5638 -3632 5702
rect -3568 5638 -3552 5702
rect -3488 5638 -3472 5702
rect -3408 5638 -3392 5702
rect -3328 5638 -3310 5702
rect -3730 5622 -3708 5638
rect -3652 5622 -3628 5638
rect -3572 5622 -3548 5638
rect -3492 5622 -3468 5638
rect -3412 5622 -3388 5638
rect -3332 5622 -3310 5638
rect -3730 5615 -3310 5622
rect -2690 5702 -2270 5720
rect -2690 5638 -2672 5702
rect -2608 5638 -2592 5702
rect -2528 5638 -2512 5702
rect -2448 5638 -2432 5702
rect -2368 5638 -2352 5702
rect -2288 5638 -2270 5702
rect -2690 5622 -2668 5638
rect -2612 5622 -2588 5638
rect -2532 5622 -2508 5638
rect -2452 5622 -2428 5638
rect -2372 5622 -2348 5638
rect -2292 5622 -2270 5638
rect -2690 5615 -2270 5622
rect -1230 5702 -810 5720
rect -1230 5638 -1212 5702
rect -1148 5638 -1132 5702
rect -1068 5638 -1052 5702
rect -988 5638 -972 5702
rect -908 5638 -892 5702
rect -828 5638 -810 5702
rect -1230 5622 -1208 5638
rect -1152 5622 -1128 5638
rect -1072 5622 -1048 5638
rect -992 5622 -968 5638
rect -912 5622 -888 5638
rect -832 5622 -810 5638
rect -1230 5615 -810 5622
rect 1810 5708 1848 5772
rect 1912 5708 1950 5772
rect 1810 5692 1950 5708
rect 1810 5628 1848 5692
rect 1912 5628 1950 5692
rect 1810 5620 1950 5628
rect -1750 4944 -1654 4950
rect -1750 4880 -1734 4944
rect -1670 4880 -1654 4944
rect -1750 4874 -1654 4880
rect -5170 4098 -4750 4105
rect -5170 4082 -5148 4098
rect -5092 4082 -5068 4098
rect -5012 4082 -4988 4098
rect -4932 4082 -4908 4098
rect -4852 4082 -4828 4098
rect -4772 4082 -4750 4098
rect -5170 4018 -5152 4082
rect -5088 4018 -5072 4082
rect -5008 4018 -4992 4082
rect -4928 4018 -4912 4082
rect -4848 4018 -4832 4082
rect -4768 4018 -4750 4082
rect -5170 4000 -4750 4018
rect -5310 3600 -5230 3605
rect -5350 3592 -5230 3600
rect -5350 3528 -5322 3592
rect -5258 3588 -5230 3592
rect -5242 3532 -5230 3588
rect -5258 3528 -5230 3532
rect -5350 3512 -5230 3528
rect -5350 3448 -5322 3512
rect -5258 3508 -5230 3512
rect -5242 3452 -5230 3508
rect -5258 3448 -5230 3452
rect -5350 3432 -5230 3448
rect -5350 3368 -5322 3432
rect -5258 3428 -5230 3432
rect -5242 3372 -5230 3428
rect -5258 3368 -5230 3372
rect -5350 3352 -5230 3368
rect -5350 3288 -5322 3352
rect -5258 3348 -5230 3352
rect -5242 3292 -5230 3348
rect -5258 3288 -5230 3292
rect -5350 3272 -5230 3288
rect -5350 3208 -5322 3272
rect -5258 3268 -5230 3272
rect -5242 3212 -5230 3268
rect -5258 3208 -5230 3212
rect -5350 3200 -5230 3208
rect -5310 3195 -5230 3200
rect -4070 3240 -3990 3245
rect -4070 3232 -3950 3240
rect -4070 3228 -4042 3232
rect -4070 3172 -4058 3228
rect -4070 3168 -4042 3172
rect -3978 3168 -3950 3232
rect -4070 3152 -3950 3168
rect -4070 3148 -4042 3152
rect -4070 3092 -4058 3148
rect -4070 3088 -4042 3092
rect -3978 3088 -3950 3152
rect -4070 3072 -3950 3088
rect -4070 3068 -4042 3072
rect -4070 3012 -4058 3068
rect -4070 3008 -4042 3012
rect -3978 3008 -3950 3072
rect -4070 2992 -3950 3008
rect -4070 2988 -4042 2992
rect -4070 2932 -4058 2988
rect -4070 2928 -4042 2932
rect -3978 2928 -3950 2992
rect -4070 2912 -3950 2928
rect -4070 2908 -4042 2912
rect -4070 2852 -4058 2908
rect -4070 2848 -4042 2852
rect -3978 2848 -3950 2912
rect -4070 2840 -3950 2848
rect -4070 2835 -3990 2840
rect -3832 2658 -3700 4300
rect -1230 4098 -810 4105
rect -1230 4082 -1208 4098
rect -1152 4082 -1128 4098
rect -1072 4082 -1048 4098
rect -992 4082 -968 4098
rect -912 4082 -888 4098
rect -832 4082 -810 4098
rect -3832 2602 -3773 2658
rect -3717 2602 -3700 2658
rect -3832 2590 -3700 2602
rect -1772 2658 -1642 4038
rect -1230 4018 -1212 4082
rect -1148 4018 -1132 4082
rect -1068 4018 -1052 4082
rect -988 4018 -972 4082
rect -908 4018 -892 4082
rect -828 4018 -810 4082
rect -1230 4000 -810 4018
rect 1810 4092 1950 4100
rect 1810 4028 1848 4092
rect 1912 4028 1950 4092
rect 1810 4012 1950 4028
rect 1810 3948 1848 4012
rect 1912 3948 1950 4012
rect 1810 3940 1950 3948
rect 1810 3920 1820 3940
rect 1940 3920 1950 3940
rect -1772 2602 -1733 2658
rect -1677 2602 -1642 2658
rect -1772 2560 -1642 2602
rect -5310 2500 -5230 2505
rect -5350 2492 -5230 2500
rect -5350 2428 -5322 2492
rect -5258 2488 -5230 2492
rect -5242 2432 -5230 2488
rect -5258 2428 -5230 2432
rect -5350 2412 -5230 2428
rect -5350 2348 -5322 2412
rect -5258 2408 -5230 2412
rect -5242 2352 -5230 2408
rect -5258 2348 -5230 2352
rect -5350 2332 -5230 2348
rect -5350 2268 -5322 2332
rect -5258 2328 -5230 2332
rect -5242 2272 -5230 2328
rect -5258 2268 -5230 2272
rect -5350 2252 -5230 2268
rect -4090 2328 -3990 2335
rect -4090 2272 -4068 2328
rect -4012 2272 -3990 2328
rect -4090 2265 -3990 2272
rect -5350 2188 -5322 2252
rect -5258 2248 -5230 2252
rect -5242 2192 -5230 2248
rect -5258 2188 -5230 2192
rect -5350 2172 -5230 2188
rect -5350 2108 -5322 2172
rect -5258 2168 -5230 2172
rect -5242 2112 -5230 2168
rect -5258 2108 -5230 2112
rect -5350 2100 -5230 2108
rect -5310 2095 -5230 2100
rect -4070 2120 -3990 2125
rect -4070 2112 -3950 2120
rect -4070 2108 -4042 2112
rect -4070 2052 -4058 2108
rect -4070 2048 -4042 2052
rect -3978 2048 -3950 2112
rect -4070 2032 -3950 2048
rect -4070 2028 -4042 2032
rect -4070 1972 -4058 2028
rect -4070 1968 -4042 1972
rect -3978 1968 -3950 2032
rect -4070 1952 -3950 1968
rect -4070 1948 -4042 1952
rect -4070 1892 -4058 1948
rect -4070 1888 -4042 1892
rect -3978 1888 -3950 1952
rect -4070 1872 -3950 1888
rect -4070 1868 -4042 1872
rect -4070 1812 -4058 1868
rect -4070 1808 -4042 1812
rect -3978 1808 -3950 1872
rect -4070 1792 -3950 1808
rect -4070 1788 -4042 1792
rect -4070 1732 -4058 1788
rect -4070 1728 -4042 1732
rect -3978 1728 -3950 1792
rect -4070 1720 -3950 1728
rect -4070 1715 -3990 1720
rect 6300 1405 6500 1800
rect 6290 1398 6510 1405
rect -5310 1380 -5230 1385
rect -5350 1372 -5230 1380
rect -5350 1308 -5322 1372
rect -5258 1368 -5230 1372
rect -5242 1312 -5230 1368
rect -5258 1308 -5230 1312
rect -5350 1292 -5230 1308
rect -5350 1228 -5322 1292
rect -5258 1288 -5230 1292
rect -5242 1232 -5230 1288
rect -5258 1228 -5230 1232
rect -5350 1212 -5230 1228
rect -5350 1148 -5322 1212
rect -5258 1208 -5230 1212
rect -5242 1152 -5230 1208
rect -5258 1148 -5230 1152
rect -5350 1132 -5230 1148
rect -5350 1068 -5322 1132
rect -5258 1128 -5230 1132
rect -5242 1072 -5230 1128
rect 6290 1102 6332 1398
rect 6468 1102 6510 1398
rect 6290 1095 6510 1102
rect -5258 1068 -5230 1072
rect -5350 1052 -5230 1068
rect -5350 988 -5322 1052
rect -5258 1048 -5230 1052
rect -5242 992 -5230 1048
rect -5258 988 -5230 992
rect -5350 980 -5230 988
rect -5310 975 -5230 980
rect -3470 822 -2750 840
rect -3470 798 -3422 822
rect -3358 798 -3342 822
rect -3278 798 -3262 822
rect -3198 798 -3182 822
rect -3118 798 -3102 822
rect -3038 798 -3022 822
rect -2958 798 -2942 822
rect -2878 798 -2862 822
rect -2798 798 -2750 822
rect -3470 742 -3458 798
rect -3402 742 -3378 758
rect -3322 742 -3298 758
rect -3242 742 -3218 758
rect -3162 742 -3138 758
rect -3082 742 -3058 758
rect -3002 742 -2978 758
rect -2922 742 -2898 758
rect -2842 742 -2818 758
rect -2762 742 -2750 798
rect -3470 735 -2750 742
rect -1080 817 -960 850
rect -1080 753 -1052 817
rect -988 753 -960 817
rect -1080 720 -960 753
rect 4810 848 5150 865
rect 4810 832 4832 848
rect 4888 832 4912 848
rect 4968 832 4992 848
rect 5048 832 5072 848
rect 5128 832 5150 848
rect 4810 768 4828 832
rect 4892 768 4908 832
rect 4972 768 4988 832
rect 5052 768 5068 832
rect 5132 768 5150 832
rect 4810 740 5150 768
<< via3 >>
rect -5152 5678 -5088 5702
rect -5152 5638 -5148 5678
rect -5148 5638 -5092 5678
rect -5092 5638 -5088 5678
rect -5072 5678 -5008 5702
rect -5072 5638 -5068 5678
rect -5068 5638 -5012 5678
rect -5012 5638 -5008 5678
rect -4992 5678 -4928 5702
rect -4992 5638 -4988 5678
rect -4988 5638 -4932 5678
rect -4932 5638 -4928 5678
rect -4912 5678 -4848 5702
rect -4912 5638 -4908 5678
rect -4908 5638 -4852 5678
rect -4852 5638 -4848 5678
rect -4832 5678 -4768 5702
rect -4832 5638 -4828 5678
rect -4828 5638 -4772 5678
rect -4772 5638 -4768 5678
rect -3712 5678 -3648 5702
rect -3712 5638 -3708 5678
rect -3708 5638 -3652 5678
rect -3652 5638 -3648 5678
rect -3632 5678 -3568 5702
rect -3632 5638 -3628 5678
rect -3628 5638 -3572 5678
rect -3572 5638 -3568 5678
rect -3552 5678 -3488 5702
rect -3552 5638 -3548 5678
rect -3548 5638 -3492 5678
rect -3492 5638 -3488 5678
rect -3472 5678 -3408 5702
rect -3472 5638 -3468 5678
rect -3468 5638 -3412 5678
rect -3412 5638 -3408 5678
rect -3392 5678 -3328 5702
rect -3392 5638 -3388 5678
rect -3388 5638 -3332 5678
rect -3332 5638 -3328 5678
rect -2672 5678 -2608 5702
rect -2672 5638 -2668 5678
rect -2668 5638 -2612 5678
rect -2612 5638 -2608 5678
rect -2592 5678 -2528 5702
rect -2592 5638 -2588 5678
rect -2588 5638 -2532 5678
rect -2532 5638 -2528 5678
rect -2512 5678 -2448 5702
rect -2512 5638 -2508 5678
rect -2508 5638 -2452 5678
rect -2452 5638 -2448 5678
rect -2432 5678 -2368 5702
rect -2432 5638 -2428 5678
rect -2428 5638 -2372 5678
rect -2372 5638 -2368 5678
rect -2352 5678 -2288 5702
rect -2352 5638 -2348 5678
rect -2348 5638 -2292 5678
rect -2292 5638 -2288 5678
rect -1212 5678 -1148 5702
rect -1212 5638 -1208 5678
rect -1208 5638 -1152 5678
rect -1152 5638 -1148 5678
rect -1132 5678 -1068 5702
rect -1132 5638 -1128 5678
rect -1128 5638 -1072 5678
rect -1072 5638 -1068 5678
rect -1052 5678 -988 5702
rect -1052 5638 -1048 5678
rect -1048 5638 -992 5678
rect -992 5638 -988 5678
rect -972 5678 -908 5702
rect -972 5638 -968 5678
rect -968 5638 -912 5678
rect -912 5638 -908 5678
rect -892 5678 -828 5702
rect -892 5638 -888 5678
rect -888 5638 -832 5678
rect -832 5638 -828 5678
rect 1848 5708 1912 5772
rect 1848 5628 1912 5692
rect -1734 4880 -1670 4944
rect -5152 4042 -5148 4082
rect -5148 4042 -5092 4082
rect -5092 4042 -5088 4082
rect -5152 4018 -5088 4042
rect -5072 4042 -5068 4082
rect -5068 4042 -5012 4082
rect -5012 4042 -5008 4082
rect -5072 4018 -5008 4042
rect -4992 4042 -4988 4082
rect -4988 4042 -4932 4082
rect -4932 4042 -4928 4082
rect -4992 4018 -4928 4042
rect -4912 4042 -4908 4082
rect -4908 4042 -4852 4082
rect -4852 4042 -4848 4082
rect -4912 4018 -4848 4042
rect -4832 4042 -4828 4082
rect -4828 4042 -4772 4082
rect -4772 4042 -4768 4082
rect -4832 4018 -4768 4042
rect -5322 3588 -5258 3592
rect -5322 3532 -5298 3588
rect -5298 3532 -5258 3588
rect -5322 3528 -5258 3532
rect -5322 3508 -5258 3512
rect -5322 3452 -5298 3508
rect -5298 3452 -5258 3508
rect -5322 3448 -5258 3452
rect -5322 3428 -5258 3432
rect -5322 3372 -5298 3428
rect -5298 3372 -5258 3428
rect -5322 3368 -5258 3372
rect -5322 3348 -5258 3352
rect -5322 3292 -5298 3348
rect -5298 3292 -5258 3348
rect -5322 3288 -5258 3292
rect -5322 3268 -5258 3272
rect -5322 3212 -5298 3268
rect -5298 3212 -5258 3268
rect -5322 3208 -5258 3212
rect -4042 3228 -3978 3232
rect -4042 3172 -4002 3228
rect -4002 3172 -3978 3228
rect -4042 3168 -3978 3172
rect -4042 3148 -3978 3152
rect -4042 3092 -4002 3148
rect -4002 3092 -3978 3148
rect -4042 3088 -3978 3092
rect -4042 3068 -3978 3072
rect -4042 3012 -4002 3068
rect -4002 3012 -3978 3068
rect -4042 3008 -3978 3012
rect -4042 2988 -3978 2992
rect -4042 2932 -4002 2988
rect -4002 2932 -3978 2988
rect -4042 2928 -3978 2932
rect -4042 2908 -3978 2912
rect -4042 2852 -4002 2908
rect -4002 2852 -3978 2908
rect -4042 2848 -3978 2852
rect -1212 4042 -1208 4082
rect -1208 4042 -1152 4082
rect -1152 4042 -1148 4082
rect -1212 4018 -1148 4042
rect -1132 4042 -1128 4082
rect -1128 4042 -1072 4082
rect -1072 4042 -1068 4082
rect -1132 4018 -1068 4042
rect -1052 4042 -1048 4082
rect -1048 4042 -992 4082
rect -992 4042 -988 4082
rect -1052 4018 -988 4042
rect -972 4042 -968 4082
rect -968 4042 -912 4082
rect -912 4042 -908 4082
rect -972 4018 -908 4042
rect -892 4042 -888 4082
rect -888 4042 -832 4082
rect -832 4042 -828 4082
rect -892 4018 -828 4042
rect 1848 4028 1912 4092
rect 1848 3948 1912 4012
rect -5322 2488 -5258 2492
rect -5322 2432 -5298 2488
rect -5298 2432 -5258 2488
rect -5322 2428 -5258 2432
rect -5322 2408 -5258 2412
rect -5322 2352 -5298 2408
rect -5298 2352 -5258 2408
rect -5322 2348 -5258 2352
rect -5322 2328 -5258 2332
rect -5322 2272 -5298 2328
rect -5298 2272 -5258 2328
rect -5322 2268 -5258 2272
rect -5322 2248 -5258 2252
rect -5322 2192 -5298 2248
rect -5298 2192 -5258 2248
rect -5322 2188 -5258 2192
rect -5322 2168 -5258 2172
rect -5322 2112 -5298 2168
rect -5298 2112 -5258 2168
rect -5322 2108 -5258 2112
rect -4042 2108 -3978 2112
rect -4042 2052 -4002 2108
rect -4002 2052 -3978 2108
rect -4042 2048 -3978 2052
rect -4042 2028 -3978 2032
rect -4042 1972 -4002 2028
rect -4002 1972 -3978 2028
rect -4042 1968 -3978 1972
rect -4042 1948 -3978 1952
rect -4042 1892 -4002 1948
rect -4002 1892 -3978 1948
rect -4042 1888 -3978 1892
rect -4042 1868 -3978 1872
rect -4042 1812 -4002 1868
rect -4002 1812 -3978 1868
rect -4042 1808 -3978 1812
rect -4042 1788 -3978 1792
rect -4042 1732 -4002 1788
rect -4002 1732 -3978 1788
rect -4042 1728 -3978 1732
rect -5322 1368 -5258 1372
rect -5322 1312 -5298 1368
rect -5298 1312 -5258 1368
rect -5322 1308 -5258 1312
rect -5322 1288 -5258 1292
rect -5322 1232 -5298 1288
rect -5298 1232 -5258 1288
rect -5322 1228 -5258 1232
rect -5322 1208 -5258 1212
rect -5322 1152 -5298 1208
rect -5298 1152 -5258 1208
rect -5322 1148 -5258 1152
rect -5322 1128 -5258 1132
rect -5322 1072 -5298 1128
rect -5298 1072 -5258 1128
rect -5322 1068 -5258 1072
rect -5322 1048 -5258 1052
rect -5322 992 -5298 1048
rect -5298 992 -5258 1048
rect -5322 988 -5258 992
rect -3422 798 -3358 822
rect -3342 798 -3278 822
rect -3262 798 -3198 822
rect -3182 798 -3118 822
rect -3102 798 -3038 822
rect -3022 798 -2958 822
rect -2942 798 -2878 822
rect -2862 798 -2798 822
rect -3422 758 -3402 798
rect -3402 758 -3378 798
rect -3378 758 -3358 798
rect -3342 758 -3322 798
rect -3322 758 -3298 798
rect -3298 758 -3278 798
rect -3262 758 -3242 798
rect -3242 758 -3218 798
rect -3218 758 -3198 798
rect -3182 758 -3162 798
rect -3162 758 -3138 798
rect -3138 758 -3118 798
rect -3102 758 -3082 798
rect -3082 758 -3058 798
rect -3058 758 -3038 798
rect -3022 758 -3002 798
rect -3002 758 -2978 798
rect -2978 758 -2958 798
rect -2942 758 -2922 798
rect -2922 758 -2898 798
rect -2898 758 -2878 798
rect -2862 758 -2842 798
rect -2842 758 -2818 798
rect -2818 758 -2798 798
rect -1052 753 -988 817
rect 4828 792 4832 832
rect 4832 792 4888 832
rect 4888 792 4892 832
rect 4828 768 4892 792
rect 4908 792 4912 832
rect 4912 792 4968 832
rect 4968 792 4972 832
rect 4908 768 4972 792
rect 4988 792 4992 832
rect 4992 792 5048 832
rect 5048 792 5052 832
rect 4988 768 5052 792
rect 5068 792 5072 832
rect 5072 792 5128 832
rect 5128 792 5132 832
rect 5068 768 5132 792
<< metal4 >>
rect -5380 5772 3000 5800
rect -5380 5708 1848 5772
rect 1912 5708 3000 5772
rect -5380 5702 3000 5708
rect -5380 5638 -5152 5702
rect -5088 5638 -5072 5702
rect -5008 5638 -4992 5702
rect -4928 5638 -4912 5702
rect -4848 5638 -4832 5702
rect -4768 5638 -3712 5702
rect -3648 5638 -3632 5702
rect -3568 5638 -3552 5702
rect -3488 5638 -3472 5702
rect -3408 5638 -3392 5702
rect -3328 5638 -2672 5702
rect -2608 5638 -2592 5702
rect -2528 5638 -2512 5702
rect -2448 5638 -2432 5702
rect -2368 5638 -2352 5702
rect -2288 5638 -1212 5702
rect -1148 5638 -1132 5702
rect -1068 5638 -1052 5702
rect -988 5638 -972 5702
rect -908 5638 -892 5702
rect -828 5692 3000 5702
rect -828 5638 1848 5692
rect -5380 5628 1848 5638
rect 1912 5628 3000 5692
rect -5380 5600 3000 5628
rect -5380 4120 -5180 5600
rect -1741 4944 -1663 4951
rect -1741 4880 -1734 4944
rect -1670 4940 -1663 4944
rect -1670 4880 3520 4940
rect -1741 4873 -1663 4880
rect -5380 4092 3000 4120
rect -5380 4082 1848 4092
rect -5380 4018 -5152 4082
rect -5088 4018 -5072 4082
rect -5008 4018 -4992 4082
rect -4928 4018 -4912 4082
rect -4848 4018 -4832 4082
rect -4768 4018 -1212 4082
rect -1148 4018 -1132 4082
rect -1068 4018 -1052 4082
rect -988 4018 -972 4082
rect -908 4018 -892 4082
rect -828 4028 1848 4082
rect 1912 4028 3000 4092
rect -828 4018 3000 4028
rect -5380 4012 3000 4018
rect -5380 3948 1848 4012
rect 1912 3948 3000 4012
rect -5380 3920 3000 3948
rect -5380 3600 3160 3800
rect -5380 3592 -5180 3600
rect -5380 3528 -5322 3592
rect -5258 3528 -5180 3592
rect -5380 3512 -5180 3528
rect -5380 3448 -5322 3512
rect -5258 3448 -5180 3512
rect -5380 3432 -5180 3448
rect -5380 3368 -5322 3432
rect -5258 3368 -5180 3432
rect -5380 3352 -5180 3368
rect -5380 3288 -5322 3352
rect -5258 3288 -5180 3352
rect -5380 3272 -5180 3288
rect -5380 3208 -5322 3272
rect -5258 3208 -5180 3272
rect -5380 2492 -5180 3208
rect -5380 2428 -5322 2492
rect -5258 2428 -5180 2492
rect -5380 2412 -5180 2428
rect -5380 2348 -5322 2412
rect -5258 2348 -5180 2412
rect -5380 2332 -5180 2348
rect -5380 2268 -5322 2332
rect -5258 2268 -5180 2332
rect -5380 2252 -5180 2268
rect -5380 2188 -5322 2252
rect -5258 2188 -5180 2252
rect -5380 2172 -5180 2188
rect -5380 2108 -5322 2172
rect -5258 2108 -5180 2172
rect -5380 1372 -5180 2108
rect -5380 1308 -5322 1372
rect -5258 1308 -5180 1372
rect -5380 1292 -5180 1308
rect -5380 1228 -5322 1292
rect -5258 1228 -5180 1292
rect -5380 1212 -5180 1228
rect -5380 1148 -5322 1212
rect -5258 1148 -5180 1212
rect -5380 1132 -5180 1148
rect -5380 1068 -5322 1132
rect -5258 1068 -5180 1132
rect -5380 1052 -5180 1068
rect -5380 988 -5322 1052
rect -5258 988 -5180 1052
rect -5380 860 -5180 988
rect -4100 3232 -3900 3600
rect -4100 3168 -4042 3232
rect -3978 3168 -3900 3232
rect -4100 3152 -3900 3168
rect -4100 3088 -4042 3152
rect -3978 3088 -3900 3152
rect -4100 3072 -3900 3088
rect -4100 3008 -4042 3072
rect -3978 3008 -3900 3072
rect -4100 2992 -3900 3008
rect -4100 2928 -4042 2992
rect -3978 2928 -3900 2992
rect -4100 2912 -3900 2928
rect -4100 2848 -4042 2912
rect -3978 2848 -3900 2912
rect -4100 2112 -3900 2848
rect -4100 2048 -4042 2112
rect -3978 2048 -3900 2112
rect -4100 2032 -3900 2048
rect -4100 1968 -4042 2032
rect -3978 1968 -3900 2032
rect -4100 1952 -3900 1968
rect -4100 1888 -4042 1952
rect -3978 1888 -3900 1952
rect -4100 1872 -3900 1888
rect -4100 1808 -4042 1872
rect -3978 1808 -3900 1872
rect -4100 1792 -3900 1808
rect -4100 1728 -4042 1792
rect -3978 1728 -3900 1792
rect -4100 860 -3900 1728
rect 4819 860 5141 861
rect -5380 832 6740 860
rect -5380 822 4828 832
rect -5380 758 -3422 822
rect -3358 758 -3342 822
rect -3278 758 -3262 822
rect -3198 758 -3182 822
rect -3118 758 -3102 822
rect -3038 758 -3022 822
rect -2958 758 -2942 822
rect -2878 758 -2862 822
rect -2798 817 4828 822
rect -2798 758 -1052 817
rect -5380 753 -1052 758
rect -988 768 4828 817
rect 4892 768 4908 832
rect 4972 768 4988 832
rect 5052 768 5068 832
rect 5132 768 6740 832
rect -988 753 6740 768
rect -5380 660 6740 753
use XM_actload2  XM_actload2_0
timestamp 1663011646
transform 1 0 -2047 0 1 753
box -43 -50 2561 3163
use XM_cs  XM_cs_0
timestamp 1663011646
transform 1 0 664 0 1 753
box -140 -53 2482 5650
use XM_diffpair  XM_diffpair_0
timestamp 1663011646
transform 1 0 -3688 0 1 2162
box -360 -1306 1506 1586
use XM_ppair  XM_ppair_0
timestamp 1663011646
transform 1 0 -5102 0 1 5030
box -220 -1060 4440 720
use XM_tail  XM_tail_0
timestamp 1663011646
transform 1 0 -5225 0 1 839
box -43 -41 1200 2921
use sky130_fd_pr__cap_mim_m3_1_EN3Q86  sky130_fd_pr__cap_mim_m3_1_EN3Q86_0
timestamp 1663011646
transform 1 0 4943 0 1 3949
box -1750 -2240 1647 2240
use sky130_fd_pr__res_high_po_2p85_7J2RPB  sky130_fd_pr__res_high_po_2p85_7J2RPB_0
timestamp 1663011646
transform 0 1 4968 -1 0 1241
box -441 -1798 441 1798
<< labels >>
rlabel metal1 s -4685 710 -750 770 4 bias_0p7
port 1 nsew
rlabel metal2 s 3009 907 3356 1047 4 out
port 2 nsew
rlabel metal2 s -2480 2590 -1740 2670 4 first_stage_out
port 3 nsew
rlabel metal3 s -3832 2660 -3700 4300 4 ppair_gate
port 4 nsew
rlabel metal4 s -820 5600 1820 5800 4 vdd
port 5 nsew
rlabel metal4 s -5380 660 -3460 860 4 vss
port 6 nsew
flabel metal2 s -2752 2172 -2652 2252 0 FreeSans 2000 0 0 0 in_n
port 7 nsew
flabel metal2 s -2752 2352 -2652 2432 0 FreeSans 2000 0 0 0 in_p
port 8 nsew
flabel metal2 s 301 2157 647 2289 0 FreeSans 2000 0 0 0 out
port 2 nsew
flabel metal1 s -1324 594 -1276 766 0 FreeSans 2000 0 0 0 bias_0p7
port 1 nsew
<< end >>
