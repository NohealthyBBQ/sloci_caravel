magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
<< pwell >>
rect -201 -300 201 300
<< nmoslvt >>
rect -15 -100 15 100
<< ndiff >>
rect -73 85 -15 100
rect -73 51 -61 85
rect -27 51 -15 85
rect -73 17 -15 51
rect -73 -17 -61 17
rect -27 -17 -15 17
rect -73 -51 -15 -17
rect -73 -85 -61 -51
rect -27 -85 -15 -51
rect -73 -100 -15 -85
rect 15 85 73 100
rect 15 51 27 85
rect 61 51 73 85
rect 15 17 73 51
rect 15 -17 27 17
rect 61 -17 73 17
rect 15 -51 73 -17
rect 15 -85 27 -51
rect 61 -85 73 -51
rect 15 -100 73 -85
<< ndiffc >>
rect -61 51 -27 85
rect -61 -17 -27 17
rect -61 -85 -27 -51
rect 27 51 61 85
rect 27 -17 61 17
rect 27 -85 61 -51
<< psubdiff >>
rect -175 240 -51 274
rect -17 240 17 274
rect 51 240 175 274
rect -175 153 -141 240
rect 141 153 175 240
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect -175 -240 -141 -153
rect 141 -240 175 -153
rect -175 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 175 -240
<< psubdiffcont >>
rect -51 240 -17 274
rect 17 240 51 274
rect -175 119 -141 153
rect 141 119 175 153
rect -175 51 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -51
rect 141 51 175 85
rect 141 -17 175 17
rect 141 -85 175 -51
rect -175 -153 -141 -119
rect 141 -153 175 -119
rect -51 -274 -17 -240
rect 17 -274 51 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -15 100 15 122
rect -15 -122 15 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -175 240 -51 274
rect -17 240 17 274
rect 51 240 175 274
rect -175 153 -141 240
rect -33 138 -17 172
rect 17 138 33 172
rect 141 153 175 240
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -61 85 -27 104
rect -61 17 -27 19
rect -61 -19 -27 -17
rect -61 -104 -27 -85
rect 27 85 61 104
rect 27 17 61 19
rect 27 -19 61 -17
rect 27 -104 61 -85
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect -175 -240 -141 -153
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect 141 -240 175 -153
rect -175 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 175 -240
<< viali >>
rect -17 138 17 172
rect -61 51 -27 53
rect -61 19 -27 51
rect -61 -51 -27 -19
rect -61 -53 -27 -51
rect 27 51 61 53
rect 27 19 61 51
rect 27 -51 61 -19
rect 27 -53 61 -51
rect -17 -172 17 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -67 53 -21 100
rect -67 19 -61 53
rect -27 19 -21 53
rect -67 -19 -21 19
rect -67 -53 -61 -19
rect -27 -53 -21 -19
rect -67 -100 -21 -53
rect 21 53 67 100
rect 21 19 27 53
rect 61 19 67 53
rect 21 -19 67 19
rect 21 -53 27 -19
rect 61 -53 67 -19
rect 21 -100 67 -53
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
<< properties >>
string FIXED_BBOX -158 -257 158 257
<< end >>
