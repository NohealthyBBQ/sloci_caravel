magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect -20 2710 130 2790
rect 1010 2710 1160 2790
rect -20 2150 130 2230
rect 1010 2150 1160 2230
rect -20 1600 130 1680
rect 1010 1590 1160 1670
rect -20 1040 130 1120
rect 1010 1040 1160 1120
rect -20 480 130 560
rect 1010 480 1160 560
<< metal1 >>
rect 530 2606 620 2610
rect 530 2554 549 2606
rect 601 2554 620 2606
rect 530 2550 620 2554
rect 330 80 370 2350
rect 537 2305 607 2351
rect 530 2056 620 2060
rect 530 2004 549 2056
rect 601 2004 620 2056
rect 530 2000 620 2004
rect 537 1749 607 1795
rect 530 1486 620 1490
rect 530 1434 549 1486
rect 601 1434 620 1486
rect 530 1430 620 1434
rect 537 1193 607 1239
rect 530 926 620 930
rect 530 874 549 926
rect 601 874 620 926
rect 530 870 620 874
rect 537 637 607 683
rect 530 386 620 390
rect 530 334 549 386
rect 601 334 620 386
rect 530 330 620 334
rect 537 81 607 127
rect 540 -40 600 81
rect 780 80 820 2350
<< via1 >>
rect 549 2554 601 2606
rect 549 2004 601 2056
rect 549 1434 601 1486
rect 549 874 601 926
rect 549 334 601 386
<< metal2 >>
rect 540 2606 610 2620
rect 540 2554 549 2606
rect 601 2554 610 2606
rect 540 2056 610 2554
rect 540 2004 549 2056
rect 601 2004 610 2056
rect 540 1500 610 2004
rect 540 1486 1200 1500
rect 540 1434 549 1486
rect 601 1434 1200 1486
rect 540 1420 1200 1434
rect 540 926 610 1420
rect 540 874 549 926
rect 601 874 610 926
rect 540 386 610 874
rect 540 334 549 386
rect 601 334 610 386
rect 540 320 610 334
use sky130_fd_pr__nfet_01v8_lvt_7MFZYU  sky130_fd_pr__nfet_01v8_lvt_7MFZYU_0
timestamp 1663011646
transform 1 0 572 0 1 1440
box -615 -1481 615 1481
<< end >>
