magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal1 >>
rect 70 736 150 740
rect 70 684 84 736
rect 136 684 150 736
rect 70 680 150 684
rect 590 736 670 740
rect 590 684 604 736
rect 656 684 670 736
rect 590 680 670 684
rect 1110 736 1190 740
rect 1110 684 1124 736
rect 1176 684 1190 736
rect 1110 680 1190 684
rect 330 576 410 580
rect 330 524 344 576
rect 396 524 410 576
rect 330 520 410 524
rect 850 576 930 580
rect 850 524 864 576
rect 916 524 930 576
rect 850 520 930 524
rect 1370 576 1450 580
rect 1370 524 1384 576
rect 1436 524 1450 576
rect 1370 520 1450 524
rect 144 448 1380 480
rect 70 376 150 380
rect 70 324 84 376
rect 136 324 150 376
rect 70 320 150 324
rect 590 376 670 380
rect 590 324 604 376
rect 656 324 670 376
rect 590 320 670 324
rect 330 216 410 220
rect 330 164 344 216
rect 396 164 410 216
rect 330 160 410 164
rect 740 119 780 448
rect 1110 376 1190 380
rect 1110 324 1124 376
rect 1176 324 1190 376
rect 1110 320 1190 324
rect 850 216 930 220
rect 850 164 864 216
rect 916 164 930 216
rect 850 160 930 164
rect 1370 216 1450 220
rect 1370 164 1384 216
rect 1436 164 1450 216
rect 1370 160 1450 164
rect 143 85 1367 119
rect 740 80 780 85
<< via1 >>
rect 84 684 136 736
rect 604 684 656 736
rect 1124 684 1176 736
rect 344 524 396 576
rect 864 524 916 576
rect 1384 524 1436 576
rect 84 324 136 376
rect 604 324 656 376
rect 344 164 396 216
rect 1124 324 1176 376
rect 864 164 916 216
rect 1384 164 1436 216
<< metal2 >>
rect 80 740 140 750
rect 600 740 660 750
rect 1120 740 1180 750
rect 80 736 1180 740
rect 80 684 84 736
rect 136 684 604 736
rect 656 684 1124 736
rect 1176 684 1180 736
rect 80 680 1180 684
rect 80 380 140 680
rect 600 670 660 680
rect 1120 670 1180 680
rect 340 580 400 590
rect 1380 580 1440 590
rect 340 576 1440 580
rect 340 524 344 576
rect 396 524 864 576
rect 916 524 1384 576
rect 1436 524 1440 576
rect 340 520 1440 524
rect 340 510 400 520
rect 600 380 660 390
rect 1120 380 1180 390
rect 80 376 1180 380
rect 80 324 84 376
rect 136 324 604 376
rect 656 324 1124 376
rect 1176 324 1180 376
rect 80 320 1180 324
rect 80 310 140 320
rect 600 310 660 320
rect 1120 310 1180 320
rect 340 220 400 230
rect 1380 220 1440 520
rect 340 216 1440 220
rect 340 164 344 216
rect 396 164 864 216
rect 916 164 1384 216
rect 1436 164 1440 216
rect 340 160 1440 164
rect 340 150 400 160
rect 1380 150 1440 160
use sky130_fd_pr__pfet_01v8_lvt_MUAP4U  sky130_fd_pr__pfet_01v8_lvt_MUAP4U_0
timestamp 1663011646
transform 1 0 759 0 1 413
box -812 -466 812 466
<< end >>
