magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -729 3542 729 3628
rect -729 -3542 -643 3542
rect 643 -3542 729 3542
rect -729 -3628 729 -3542
<< psubdiff >>
rect -703 3568 -595 3602
rect -561 3568 -527 3602
rect -493 3568 -459 3602
rect -425 3568 -391 3602
rect -357 3568 -323 3602
rect -289 3568 -255 3602
rect -221 3568 -187 3602
rect -153 3568 -119 3602
rect -85 3568 -51 3602
rect -17 3568 17 3602
rect 51 3568 85 3602
rect 119 3568 153 3602
rect 187 3568 221 3602
rect 255 3568 289 3602
rect 323 3568 357 3602
rect 391 3568 425 3602
rect 459 3568 493 3602
rect 527 3568 561 3602
rect 595 3568 703 3602
rect -703 3485 -669 3568
rect 669 3485 703 3568
rect -703 3417 -669 3451
rect -703 3349 -669 3383
rect -703 3281 -669 3315
rect -703 3213 -669 3247
rect -703 3145 -669 3179
rect -703 3077 -669 3111
rect -703 3009 -669 3043
rect -703 2941 -669 2975
rect -703 2873 -669 2907
rect -703 2805 -669 2839
rect -703 2737 -669 2771
rect -703 2669 -669 2703
rect -703 2601 -669 2635
rect -703 2533 -669 2567
rect -703 2465 -669 2499
rect -703 2397 -669 2431
rect -703 2329 -669 2363
rect -703 2261 -669 2295
rect -703 2193 -669 2227
rect -703 2125 -669 2159
rect -703 2057 -669 2091
rect -703 1989 -669 2023
rect -703 1921 -669 1955
rect -703 1853 -669 1887
rect -703 1785 -669 1819
rect -703 1717 -669 1751
rect -703 1649 -669 1683
rect -703 1581 -669 1615
rect -703 1513 -669 1547
rect -703 1445 -669 1479
rect -703 1377 -669 1411
rect -703 1309 -669 1343
rect -703 1241 -669 1275
rect -703 1173 -669 1207
rect -703 1105 -669 1139
rect -703 1037 -669 1071
rect -703 969 -669 1003
rect -703 901 -669 935
rect -703 833 -669 867
rect -703 765 -669 799
rect -703 697 -669 731
rect -703 629 -669 663
rect -703 561 -669 595
rect -703 493 -669 527
rect -703 425 -669 459
rect -703 357 -669 391
rect -703 289 -669 323
rect -703 221 -669 255
rect -703 153 -669 187
rect -703 85 -669 119
rect -703 17 -669 51
rect -703 -51 -669 -17
rect -703 -119 -669 -85
rect -703 -187 -669 -153
rect -703 -255 -669 -221
rect -703 -323 -669 -289
rect -703 -391 -669 -357
rect -703 -459 -669 -425
rect -703 -527 -669 -493
rect -703 -595 -669 -561
rect -703 -663 -669 -629
rect -703 -731 -669 -697
rect -703 -799 -669 -765
rect -703 -867 -669 -833
rect -703 -935 -669 -901
rect -703 -1003 -669 -969
rect -703 -1071 -669 -1037
rect -703 -1139 -669 -1105
rect -703 -1207 -669 -1173
rect -703 -1275 -669 -1241
rect -703 -1343 -669 -1309
rect -703 -1411 -669 -1377
rect -703 -1479 -669 -1445
rect -703 -1547 -669 -1513
rect -703 -1615 -669 -1581
rect -703 -1683 -669 -1649
rect -703 -1751 -669 -1717
rect -703 -1819 -669 -1785
rect -703 -1887 -669 -1853
rect -703 -1955 -669 -1921
rect -703 -2023 -669 -1989
rect -703 -2091 -669 -2057
rect -703 -2159 -669 -2125
rect -703 -2227 -669 -2193
rect -703 -2295 -669 -2261
rect -703 -2363 -669 -2329
rect -703 -2431 -669 -2397
rect -703 -2499 -669 -2465
rect -703 -2567 -669 -2533
rect -703 -2635 -669 -2601
rect -703 -2703 -669 -2669
rect -703 -2771 -669 -2737
rect -703 -2839 -669 -2805
rect -703 -2907 -669 -2873
rect -703 -2975 -669 -2941
rect -703 -3043 -669 -3009
rect -703 -3111 -669 -3077
rect -703 -3179 -669 -3145
rect -703 -3247 -669 -3213
rect -703 -3315 -669 -3281
rect -703 -3383 -669 -3349
rect -703 -3451 -669 -3417
rect 669 3417 703 3451
rect 669 3349 703 3383
rect 669 3281 703 3315
rect 669 3213 703 3247
rect 669 3145 703 3179
rect 669 3077 703 3111
rect 669 3009 703 3043
rect 669 2941 703 2975
rect 669 2873 703 2907
rect 669 2805 703 2839
rect 669 2737 703 2771
rect 669 2669 703 2703
rect 669 2601 703 2635
rect 669 2533 703 2567
rect 669 2465 703 2499
rect 669 2397 703 2431
rect 669 2329 703 2363
rect 669 2261 703 2295
rect 669 2193 703 2227
rect 669 2125 703 2159
rect 669 2057 703 2091
rect 669 1989 703 2023
rect 669 1921 703 1955
rect 669 1853 703 1887
rect 669 1785 703 1819
rect 669 1717 703 1751
rect 669 1649 703 1683
rect 669 1581 703 1615
rect 669 1513 703 1547
rect 669 1445 703 1479
rect 669 1377 703 1411
rect 669 1309 703 1343
rect 669 1241 703 1275
rect 669 1173 703 1207
rect 669 1105 703 1139
rect 669 1037 703 1071
rect 669 969 703 1003
rect 669 901 703 935
rect 669 833 703 867
rect 669 765 703 799
rect 669 697 703 731
rect 669 629 703 663
rect 669 561 703 595
rect 669 493 703 527
rect 669 425 703 459
rect 669 357 703 391
rect 669 289 703 323
rect 669 221 703 255
rect 669 153 703 187
rect 669 85 703 119
rect 669 17 703 51
rect 669 -51 703 -17
rect 669 -119 703 -85
rect 669 -187 703 -153
rect 669 -255 703 -221
rect 669 -323 703 -289
rect 669 -391 703 -357
rect 669 -459 703 -425
rect 669 -527 703 -493
rect 669 -595 703 -561
rect 669 -663 703 -629
rect 669 -731 703 -697
rect 669 -799 703 -765
rect 669 -867 703 -833
rect 669 -935 703 -901
rect 669 -1003 703 -969
rect 669 -1071 703 -1037
rect 669 -1139 703 -1105
rect 669 -1207 703 -1173
rect 669 -1275 703 -1241
rect 669 -1343 703 -1309
rect 669 -1411 703 -1377
rect 669 -1479 703 -1445
rect 669 -1547 703 -1513
rect 669 -1615 703 -1581
rect 669 -1683 703 -1649
rect 669 -1751 703 -1717
rect 669 -1819 703 -1785
rect 669 -1887 703 -1853
rect 669 -1955 703 -1921
rect 669 -2023 703 -1989
rect 669 -2091 703 -2057
rect 669 -2159 703 -2125
rect 669 -2227 703 -2193
rect 669 -2295 703 -2261
rect 669 -2363 703 -2329
rect 669 -2431 703 -2397
rect 669 -2499 703 -2465
rect 669 -2567 703 -2533
rect 669 -2635 703 -2601
rect 669 -2703 703 -2669
rect 669 -2771 703 -2737
rect 669 -2839 703 -2805
rect 669 -2907 703 -2873
rect 669 -2975 703 -2941
rect 669 -3043 703 -3009
rect 669 -3111 703 -3077
rect 669 -3179 703 -3145
rect 669 -3247 703 -3213
rect 669 -3315 703 -3281
rect 669 -3383 703 -3349
rect 669 -3451 703 -3417
rect -703 -3568 -669 -3485
rect 669 -3568 703 -3485
rect -703 -3602 -595 -3568
rect -561 -3602 -527 -3568
rect -493 -3602 -459 -3568
rect -425 -3602 -391 -3568
rect -357 -3602 -323 -3568
rect -289 -3602 -255 -3568
rect -221 -3602 -187 -3568
rect -153 -3602 -119 -3568
rect -85 -3602 -51 -3568
rect -17 -3602 17 -3568
rect 51 -3602 85 -3568
rect 119 -3602 153 -3568
rect 187 -3602 221 -3568
rect 255 -3602 289 -3568
rect 323 -3602 357 -3568
rect 391 -3602 425 -3568
rect 459 -3602 493 -3568
rect 527 -3602 561 -3568
rect 595 -3602 703 -3568
<< psubdiffcont >>
rect -595 3568 -561 3602
rect -527 3568 -493 3602
rect -459 3568 -425 3602
rect -391 3568 -357 3602
rect -323 3568 -289 3602
rect -255 3568 -221 3602
rect -187 3568 -153 3602
rect -119 3568 -85 3602
rect -51 3568 -17 3602
rect 17 3568 51 3602
rect 85 3568 119 3602
rect 153 3568 187 3602
rect 221 3568 255 3602
rect 289 3568 323 3602
rect 357 3568 391 3602
rect 425 3568 459 3602
rect 493 3568 527 3602
rect 561 3568 595 3602
rect -703 3451 -669 3485
rect -703 3383 -669 3417
rect -703 3315 -669 3349
rect -703 3247 -669 3281
rect -703 3179 -669 3213
rect -703 3111 -669 3145
rect -703 3043 -669 3077
rect -703 2975 -669 3009
rect -703 2907 -669 2941
rect -703 2839 -669 2873
rect -703 2771 -669 2805
rect -703 2703 -669 2737
rect -703 2635 -669 2669
rect -703 2567 -669 2601
rect -703 2499 -669 2533
rect -703 2431 -669 2465
rect -703 2363 -669 2397
rect -703 2295 -669 2329
rect -703 2227 -669 2261
rect -703 2159 -669 2193
rect -703 2091 -669 2125
rect -703 2023 -669 2057
rect -703 1955 -669 1989
rect -703 1887 -669 1921
rect -703 1819 -669 1853
rect -703 1751 -669 1785
rect -703 1683 -669 1717
rect -703 1615 -669 1649
rect -703 1547 -669 1581
rect -703 1479 -669 1513
rect -703 1411 -669 1445
rect -703 1343 -669 1377
rect -703 1275 -669 1309
rect -703 1207 -669 1241
rect -703 1139 -669 1173
rect -703 1071 -669 1105
rect -703 1003 -669 1037
rect -703 935 -669 969
rect -703 867 -669 901
rect -703 799 -669 833
rect -703 731 -669 765
rect -703 663 -669 697
rect -703 595 -669 629
rect -703 527 -669 561
rect -703 459 -669 493
rect -703 391 -669 425
rect -703 323 -669 357
rect -703 255 -669 289
rect -703 187 -669 221
rect -703 119 -669 153
rect -703 51 -669 85
rect -703 -17 -669 17
rect -703 -85 -669 -51
rect -703 -153 -669 -119
rect -703 -221 -669 -187
rect -703 -289 -669 -255
rect -703 -357 -669 -323
rect -703 -425 -669 -391
rect -703 -493 -669 -459
rect -703 -561 -669 -527
rect -703 -629 -669 -595
rect -703 -697 -669 -663
rect -703 -765 -669 -731
rect -703 -833 -669 -799
rect -703 -901 -669 -867
rect -703 -969 -669 -935
rect -703 -1037 -669 -1003
rect -703 -1105 -669 -1071
rect -703 -1173 -669 -1139
rect -703 -1241 -669 -1207
rect -703 -1309 -669 -1275
rect -703 -1377 -669 -1343
rect -703 -1445 -669 -1411
rect -703 -1513 -669 -1479
rect -703 -1581 -669 -1547
rect -703 -1649 -669 -1615
rect -703 -1717 -669 -1683
rect -703 -1785 -669 -1751
rect -703 -1853 -669 -1819
rect -703 -1921 -669 -1887
rect -703 -1989 -669 -1955
rect -703 -2057 -669 -2023
rect -703 -2125 -669 -2091
rect -703 -2193 -669 -2159
rect -703 -2261 -669 -2227
rect -703 -2329 -669 -2295
rect -703 -2397 -669 -2363
rect -703 -2465 -669 -2431
rect -703 -2533 -669 -2499
rect -703 -2601 -669 -2567
rect -703 -2669 -669 -2635
rect -703 -2737 -669 -2703
rect -703 -2805 -669 -2771
rect -703 -2873 -669 -2839
rect -703 -2941 -669 -2907
rect -703 -3009 -669 -2975
rect -703 -3077 -669 -3043
rect -703 -3145 -669 -3111
rect -703 -3213 -669 -3179
rect -703 -3281 -669 -3247
rect -703 -3349 -669 -3315
rect -703 -3417 -669 -3383
rect -703 -3485 -669 -3451
rect 669 3451 703 3485
rect 669 3383 703 3417
rect 669 3315 703 3349
rect 669 3247 703 3281
rect 669 3179 703 3213
rect 669 3111 703 3145
rect 669 3043 703 3077
rect 669 2975 703 3009
rect 669 2907 703 2941
rect 669 2839 703 2873
rect 669 2771 703 2805
rect 669 2703 703 2737
rect 669 2635 703 2669
rect 669 2567 703 2601
rect 669 2499 703 2533
rect 669 2431 703 2465
rect 669 2363 703 2397
rect 669 2295 703 2329
rect 669 2227 703 2261
rect 669 2159 703 2193
rect 669 2091 703 2125
rect 669 2023 703 2057
rect 669 1955 703 1989
rect 669 1887 703 1921
rect 669 1819 703 1853
rect 669 1751 703 1785
rect 669 1683 703 1717
rect 669 1615 703 1649
rect 669 1547 703 1581
rect 669 1479 703 1513
rect 669 1411 703 1445
rect 669 1343 703 1377
rect 669 1275 703 1309
rect 669 1207 703 1241
rect 669 1139 703 1173
rect 669 1071 703 1105
rect 669 1003 703 1037
rect 669 935 703 969
rect 669 867 703 901
rect 669 799 703 833
rect 669 731 703 765
rect 669 663 703 697
rect 669 595 703 629
rect 669 527 703 561
rect 669 459 703 493
rect 669 391 703 425
rect 669 323 703 357
rect 669 255 703 289
rect 669 187 703 221
rect 669 119 703 153
rect 669 51 703 85
rect 669 -17 703 17
rect 669 -85 703 -51
rect 669 -153 703 -119
rect 669 -221 703 -187
rect 669 -289 703 -255
rect 669 -357 703 -323
rect 669 -425 703 -391
rect 669 -493 703 -459
rect 669 -561 703 -527
rect 669 -629 703 -595
rect 669 -697 703 -663
rect 669 -765 703 -731
rect 669 -833 703 -799
rect 669 -901 703 -867
rect 669 -969 703 -935
rect 669 -1037 703 -1003
rect 669 -1105 703 -1071
rect 669 -1173 703 -1139
rect 669 -1241 703 -1207
rect 669 -1309 703 -1275
rect 669 -1377 703 -1343
rect 669 -1445 703 -1411
rect 669 -1513 703 -1479
rect 669 -1581 703 -1547
rect 669 -1649 703 -1615
rect 669 -1717 703 -1683
rect 669 -1785 703 -1751
rect 669 -1853 703 -1819
rect 669 -1921 703 -1887
rect 669 -1989 703 -1955
rect 669 -2057 703 -2023
rect 669 -2125 703 -2091
rect 669 -2193 703 -2159
rect 669 -2261 703 -2227
rect 669 -2329 703 -2295
rect 669 -2397 703 -2363
rect 669 -2465 703 -2431
rect 669 -2533 703 -2499
rect 669 -2601 703 -2567
rect 669 -2669 703 -2635
rect 669 -2737 703 -2703
rect 669 -2805 703 -2771
rect 669 -2873 703 -2839
rect 669 -2941 703 -2907
rect 669 -3009 703 -2975
rect 669 -3077 703 -3043
rect 669 -3145 703 -3111
rect 669 -3213 703 -3179
rect 669 -3281 703 -3247
rect 669 -3349 703 -3315
rect 669 -3417 703 -3383
rect 669 -3485 703 -3451
rect -595 -3602 -561 -3568
rect -527 -3602 -493 -3568
rect -459 -3602 -425 -3568
rect -391 -3602 -357 -3568
rect -323 -3602 -289 -3568
rect -255 -3602 -221 -3568
rect -187 -3602 -153 -3568
rect -119 -3602 -85 -3568
rect -51 -3602 -17 -3568
rect 17 -3602 51 -3568
rect 85 -3602 119 -3568
rect 153 -3602 187 -3568
rect 221 -3602 255 -3568
rect 289 -3602 323 -3568
rect 357 -3602 391 -3568
rect 425 -3602 459 -3568
rect 493 -3602 527 -3568
rect 561 -3602 595 -3568
<< xpolycontact >>
rect -573 3040 573 3472
rect -573 -3472 573 -3040
<< ppolyres >>
rect -573 -3040 573 3040
<< locali >>
rect -703 3568 -595 3602
rect -561 3568 -527 3602
rect -493 3568 -459 3602
rect -425 3568 -391 3602
rect -357 3568 -323 3602
rect -289 3568 -255 3602
rect -221 3568 -187 3602
rect -153 3568 -119 3602
rect -85 3568 -51 3602
rect -17 3568 17 3602
rect 51 3568 85 3602
rect 119 3568 153 3602
rect 187 3568 221 3602
rect 255 3568 289 3602
rect 323 3568 357 3602
rect 391 3568 425 3602
rect 459 3568 493 3602
rect 527 3568 561 3602
rect 595 3568 703 3602
rect -703 3485 -669 3568
rect 669 3485 703 3568
rect -703 3417 -669 3451
rect -703 3349 -669 3383
rect -703 3281 -669 3315
rect -703 3213 -669 3247
rect -703 3145 -669 3179
rect -703 3077 -669 3111
rect -703 3009 -669 3043
rect 669 3417 703 3451
rect 669 3349 703 3383
rect 669 3281 703 3315
rect 669 3213 703 3247
rect 669 3145 703 3179
rect 669 3077 703 3111
rect -703 2941 -669 2975
rect -703 2873 -669 2907
rect -703 2805 -669 2839
rect -703 2737 -669 2771
rect -703 2669 -669 2703
rect -703 2601 -669 2635
rect -703 2533 -669 2567
rect -703 2465 -669 2499
rect -703 2397 -669 2431
rect -703 2329 -669 2363
rect -703 2261 -669 2295
rect -703 2193 -669 2227
rect -703 2125 -669 2159
rect -703 2057 -669 2091
rect -703 1989 -669 2023
rect -703 1921 -669 1955
rect -703 1853 -669 1887
rect -703 1785 -669 1819
rect -703 1717 -669 1751
rect -703 1649 -669 1683
rect -703 1581 -669 1615
rect -703 1513 -669 1547
rect -703 1445 -669 1479
rect -703 1377 -669 1411
rect -703 1309 -669 1343
rect -703 1241 -669 1275
rect -703 1173 -669 1207
rect -703 1105 -669 1139
rect -703 1037 -669 1071
rect -703 969 -669 1003
rect -703 901 -669 935
rect -703 833 -669 867
rect -703 765 -669 799
rect -703 697 -669 731
rect -703 629 -669 663
rect -703 561 -669 595
rect -703 493 -669 527
rect -703 425 -669 459
rect -703 357 -669 391
rect -703 289 -669 323
rect -703 221 -669 255
rect -703 153 -669 187
rect -703 85 -669 119
rect -703 17 -669 51
rect -703 -51 -669 -17
rect -703 -119 -669 -85
rect -703 -187 -669 -153
rect -703 -255 -669 -221
rect -703 -323 -669 -289
rect -703 -391 -669 -357
rect -703 -459 -669 -425
rect -703 -527 -669 -493
rect -703 -595 -669 -561
rect -703 -663 -669 -629
rect -703 -731 -669 -697
rect -703 -799 -669 -765
rect -703 -867 -669 -833
rect -703 -935 -669 -901
rect -703 -1003 -669 -969
rect -703 -1071 -669 -1037
rect -703 -1139 -669 -1105
rect -703 -1207 -669 -1173
rect -703 -1275 -669 -1241
rect -703 -1343 -669 -1309
rect -703 -1411 -669 -1377
rect -703 -1479 -669 -1445
rect -703 -1547 -669 -1513
rect -703 -1615 -669 -1581
rect -703 -1683 -669 -1649
rect -703 -1751 -669 -1717
rect -703 -1819 -669 -1785
rect -703 -1887 -669 -1853
rect -703 -1955 -669 -1921
rect -703 -2023 -669 -1989
rect -703 -2091 -669 -2057
rect -703 -2159 -669 -2125
rect -703 -2227 -669 -2193
rect -703 -2295 -669 -2261
rect -703 -2363 -669 -2329
rect -703 -2431 -669 -2397
rect -703 -2499 -669 -2465
rect -703 -2567 -669 -2533
rect -703 -2635 -669 -2601
rect -703 -2703 -669 -2669
rect -703 -2771 -669 -2737
rect -703 -2839 -669 -2805
rect -703 -2907 -669 -2873
rect -703 -2975 -669 -2941
rect -703 -3043 -669 -3009
rect 669 3009 703 3043
rect 669 2941 703 2975
rect 669 2873 703 2907
rect 669 2805 703 2839
rect 669 2737 703 2771
rect 669 2669 703 2703
rect 669 2601 703 2635
rect 669 2533 703 2567
rect 669 2465 703 2499
rect 669 2397 703 2431
rect 669 2329 703 2363
rect 669 2261 703 2295
rect 669 2193 703 2227
rect 669 2125 703 2159
rect 669 2057 703 2091
rect 669 1989 703 2023
rect 669 1921 703 1955
rect 669 1853 703 1887
rect 669 1785 703 1819
rect 669 1717 703 1751
rect 669 1649 703 1683
rect 669 1581 703 1615
rect 669 1513 703 1547
rect 669 1445 703 1479
rect 669 1377 703 1411
rect 669 1309 703 1343
rect 669 1241 703 1275
rect 669 1173 703 1207
rect 669 1105 703 1139
rect 669 1037 703 1071
rect 669 969 703 1003
rect 669 901 703 935
rect 669 833 703 867
rect 669 765 703 799
rect 669 697 703 731
rect 669 629 703 663
rect 669 561 703 595
rect 669 493 703 527
rect 669 425 703 459
rect 669 357 703 391
rect 669 289 703 323
rect 669 221 703 255
rect 669 153 703 187
rect 669 85 703 119
rect 669 17 703 51
rect 669 -51 703 -17
rect 669 -119 703 -85
rect 669 -187 703 -153
rect 669 -255 703 -221
rect 669 -323 703 -289
rect 669 -391 703 -357
rect 669 -459 703 -425
rect 669 -527 703 -493
rect 669 -595 703 -561
rect 669 -663 703 -629
rect 669 -731 703 -697
rect 669 -799 703 -765
rect 669 -867 703 -833
rect 669 -935 703 -901
rect 669 -1003 703 -969
rect 669 -1071 703 -1037
rect 669 -1139 703 -1105
rect 669 -1207 703 -1173
rect 669 -1275 703 -1241
rect 669 -1343 703 -1309
rect 669 -1411 703 -1377
rect 669 -1479 703 -1445
rect 669 -1547 703 -1513
rect 669 -1615 703 -1581
rect 669 -1683 703 -1649
rect 669 -1751 703 -1717
rect 669 -1819 703 -1785
rect 669 -1887 703 -1853
rect 669 -1955 703 -1921
rect 669 -2023 703 -1989
rect 669 -2091 703 -2057
rect 669 -2159 703 -2125
rect 669 -2227 703 -2193
rect 669 -2295 703 -2261
rect 669 -2363 703 -2329
rect 669 -2431 703 -2397
rect 669 -2499 703 -2465
rect 669 -2567 703 -2533
rect 669 -2635 703 -2601
rect 669 -2703 703 -2669
rect 669 -2771 703 -2737
rect 669 -2839 703 -2805
rect 669 -2907 703 -2873
rect 669 -2975 703 -2941
rect -703 -3111 -669 -3077
rect -703 -3179 -669 -3145
rect -703 -3247 -669 -3213
rect -703 -3315 -669 -3281
rect -703 -3383 -669 -3349
rect -703 -3451 -669 -3417
rect 669 -3043 703 -3009
rect 669 -3111 703 -3077
rect 669 -3179 703 -3145
rect 669 -3247 703 -3213
rect 669 -3315 703 -3281
rect 669 -3383 703 -3349
rect 669 -3451 703 -3417
rect -703 -3568 -669 -3485
rect 669 -3568 703 -3485
rect -703 -3602 -595 -3568
rect -561 -3602 -527 -3568
rect -493 -3602 -459 -3568
rect -425 -3602 -391 -3568
rect -357 -3602 -323 -3568
rect -289 -3602 -255 -3568
rect -221 -3602 -187 -3568
rect -153 -3602 -119 -3568
rect -85 -3602 -51 -3568
rect -17 -3602 17 -3568
rect 51 -3602 85 -3568
rect 119 -3602 153 -3568
rect 187 -3602 221 -3568
rect 255 -3602 289 -3568
rect 323 -3602 357 -3568
rect 391 -3602 425 -3568
rect 459 -3602 493 -3568
rect 527 -3602 561 -3568
rect 595 -3602 703 -3568
<< viali >>
rect -557 3058 557 3452
rect -557 -3453 557 -3059
<< metal1 >>
rect -569 3452 569 3460
rect -569 3058 -557 3452
rect 557 3058 569 3452
rect -569 3051 569 3058
rect -569 -3059 569 -3051
rect -569 -3453 -557 -3059
rect 557 -3453 569 -3059
rect -569 -3460 569 -3453
<< properties >>
string FIXED_BBOX -686 -3585 686 3585
<< end >>
