magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -365 172 -307 178
rect -173 172 -115 178
rect 19 172 77 178
rect 211 172 269 178
rect 403 172 461 178
rect -365 138 -353 172
rect -173 138 -161 172
rect 19 138 31 172
rect 211 138 223 172
rect 403 138 415 172
rect -365 132 -307 138
rect -173 132 -115 138
rect 19 132 77 138
rect 211 132 269 138
rect 403 132 461 138
rect -461 -138 -403 -132
rect -269 -138 -211 -132
rect -77 -138 -19 -132
rect 115 -138 173 -132
rect 307 -138 365 -132
rect -461 -172 -449 -138
rect -269 -172 -257 -138
rect -77 -172 -65 -138
rect 115 -172 127 -138
rect 307 -172 319 -138
rect -461 -178 -403 -172
rect -269 -178 -211 -172
rect -77 -178 -19 -172
rect 115 -178 173 -172
rect 307 -178 365 -172
<< pwell >>
rect -637 -300 637 300
<< nmoslvt >>
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
<< ndiff >>
rect -509 85 -447 100
rect -509 51 -497 85
rect -463 51 -447 85
rect -509 17 -447 51
rect -509 -17 -497 17
rect -463 -17 -447 17
rect -509 -51 -447 -17
rect -509 -85 -497 -51
rect -463 -85 -447 -51
rect -509 -100 -447 -85
rect -417 85 -351 100
rect -417 51 -401 85
rect -367 51 -351 85
rect -417 17 -351 51
rect -417 -17 -401 17
rect -367 -17 -351 17
rect -417 -51 -351 -17
rect -417 -85 -401 -51
rect -367 -85 -351 -51
rect -417 -100 -351 -85
rect -321 85 -255 100
rect -321 51 -305 85
rect -271 51 -255 85
rect -321 17 -255 51
rect -321 -17 -305 17
rect -271 -17 -255 17
rect -321 -51 -255 -17
rect -321 -85 -305 -51
rect -271 -85 -255 -51
rect -321 -100 -255 -85
rect -225 85 -159 100
rect -225 51 -209 85
rect -175 51 -159 85
rect -225 17 -159 51
rect -225 -17 -209 17
rect -175 -17 -159 17
rect -225 -51 -159 -17
rect -225 -85 -209 -51
rect -175 -85 -159 -51
rect -225 -100 -159 -85
rect -129 85 -63 100
rect -129 51 -113 85
rect -79 51 -63 85
rect -129 17 -63 51
rect -129 -17 -113 17
rect -79 -17 -63 17
rect -129 -51 -63 -17
rect -129 -85 -113 -51
rect -79 -85 -63 -51
rect -129 -100 -63 -85
rect -33 85 33 100
rect -33 51 -17 85
rect 17 51 33 85
rect -33 17 33 51
rect -33 -17 -17 17
rect 17 -17 33 17
rect -33 -51 33 -17
rect -33 -85 -17 -51
rect 17 -85 33 -51
rect -33 -100 33 -85
rect 63 85 129 100
rect 63 51 79 85
rect 113 51 129 85
rect 63 17 129 51
rect 63 -17 79 17
rect 113 -17 129 17
rect 63 -51 129 -17
rect 63 -85 79 -51
rect 113 -85 129 -51
rect 63 -100 129 -85
rect 159 85 225 100
rect 159 51 175 85
rect 209 51 225 85
rect 159 17 225 51
rect 159 -17 175 17
rect 209 -17 225 17
rect 159 -51 225 -17
rect 159 -85 175 -51
rect 209 -85 225 -51
rect 159 -100 225 -85
rect 255 85 321 100
rect 255 51 271 85
rect 305 51 321 85
rect 255 17 321 51
rect 255 -17 271 17
rect 305 -17 321 17
rect 255 -51 321 -17
rect 255 -85 271 -51
rect 305 -85 321 -51
rect 255 -100 321 -85
rect 351 85 417 100
rect 351 51 367 85
rect 401 51 417 85
rect 351 17 417 51
rect 351 -17 367 17
rect 401 -17 417 17
rect 351 -51 417 -17
rect 351 -85 367 -51
rect 401 -85 417 -51
rect 351 -100 417 -85
rect 447 85 509 100
rect 447 51 463 85
rect 497 51 509 85
rect 447 17 509 51
rect 447 -17 463 17
rect 497 -17 509 17
rect 447 -51 509 -17
rect 447 -85 463 -51
rect 497 -85 509 -51
rect 447 -100 509 -85
<< ndiffc >>
rect -497 51 -463 85
rect -497 -17 -463 17
rect -497 -85 -463 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -305 51 -271 85
rect -305 -17 -271 17
rect -305 -85 -271 -51
rect -209 51 -175 85
rect -209 -17 -175 17
rect -209 -85 -175 -51
rect -113 51 -79 85
rect -113 -17 -79 17
rect -113 -85 -79 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 79 51 113 85
rect 79 -17 113 17
rect 79 -85 113 -51
rect 175 51 209 85
rect 175 -17 209 17
rect 175 -85 209 -51
rect 271 51 305 85
rect 271 -17 305 17
rect 271 -85 305 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 463 51 497 85
rect 463 -17 497 17
rect 463 -85 497 -51
<< psubdiff >>
rect -611 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 611 274
rect -611 153 -577 240
rect -611 85 -577 119
rect 577 153 611 240
rect -611 17 -577 51
rect -611 -51 -577 -17
rect -611 -119 -577 -85
rect 577 85 611 119
rect 577 17 611 51
rect 577 -51 611 -17
rect -611 -240 -577 -153
rect 577 -119 611 -85
rect 577 -240 611 -153
rect -611 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 611 -240
<< psubdiffcont >>
rect -493 240 -459 274
rect -425 240 -391 274
rect -357 240 -323 274
rect -289 240 -255 274
rect -221 240 -187 274
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect 187 240 221 274
rect 255 240 289 274
rect 323 240 357 274
rect 391 240 425 274
rect 459 240 493 274
rect -611 119 -577 153
rect 577 119 611 153
rect -611 51 -577 85
rect -611 -17 -577 17
rect -611 -85 -577 -51
rect 577 51 611 85
rect 577 -17 611 17
rect 577 -85 611 -51
rect -611 -153 -577 -119
rect 577 -153 611 -119
rect -493 -274 -459 -240
rect -425 -274 -391 -240
rect -357 -274 -323 -240
rect -289 -274 -255 -240
rect -221 -274 -187 -240
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
rect 187 -274 221 -240
rect 255 -274 289 -240
rect 323 -274 357 -240
rect 391 -274 425 -240
rect 459 -274 493 -240
<< poly >>
rect -369 172 -303 188
rect -369 138 -353 172
rect -319 138 -303 172
rect -447 100 -417 126
rect -369 122 -303 138
rect -177 172 -111 188
rect -177 138 -161 172
rect -127 138 -111 172
rect -351 100 -321 122
rect -255 100 -225 126
rect -177 122 -111 138
rect 15 172 81 188
rect 15 138 31 172
rect 65 138 81 172
rect -159 100 -129 122
rect -63 100 -33 126
rect 15 122 81 138
rect 207 172 273 188
rect 207 138 223 172
rect 257 138 273 172
rect 33 100 63 122
rect 129 100 159 126
rect 207 122 273 138
rect 399 172 465 188
rect 399 138 415 172
rect 449 138 465 172
rect 225 100 255 122
rect 321 100 351 126
rect 399 122 465 138
rect 417 100 447 122
rect -447 -122 -417 -100
rect -465 -138 -399 -122
rect -351 -126 -321 -100
rect -255 -122 -225 -100
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -465 -188 -399 -172
rect -273 -138 -207 -122
rect -159 -126 -129 -100
rect -63 -122 -33 -100
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -273 -188 -207 -172
rect -81 -138 -15 -122
rect 33 -126 63 -100
rect 129 -122 159 -100
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect -81 -188 -15 -172
rect 111 -138 177 -122
rect 225 -126 255 -100
rect 321 -122 351 -100
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 111 -188 177 -172
rect 303 -138 369 -122
rect 417 -126 447 -100
rect 303 -172 319 -138
rect 353 -172 369 -138
rect 303 -188 369 -172
<< polycont >>
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
<< locali >>
rect -611 240 -493 274
rect -459 240 -425 274
rect -391 240 -357 274
rect -323 240 -289 274
rect -255 240 -221 274
rect -187 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 187 274
rect 221 240 255 274
rect 289 240 323 274
rect 357 240 391 274
rect 425 240 459 274
rect 493 240 611 274
rect -611 153 -577 240
rect -369 138 -353 172
rect -319 138 -303 172
rect -177 138 -161 172
rect -127 138 -111 172
rect 15 138 31 172
rect 65 138 81 172
rect 207 138 223 172
rect 257 138 273 172
rect 399 138 415 172
rect 449 138 465 172
rect 577 153 611 240
rect -611 85 -577 119
rect -611 17 -577 51
rect -611 -51 -577 -17
rect -611 -119 -577 -85
rect -497 85 -463 104
rect -497 17 -463 19
rect -497 -19 -463 -17
rect -497 -104 -463 -85
rect -401 85 -367 104
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -104 -367 -85
rect -305 85 -271 104
rect -305 17 -271 19
rect -305 -19 -271 -17
rect -305 -104 -271 -85
rect -209 85 -175 104
rect -209 17 -175 19
rect -209 -19 -175 -17
rect -209 -104 -175 -85
rect -113 85 -79 104
rect -113 17 -79 19
rect -113 -19 -79 -17
rect -113 -104 -79 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 79 85 113 104
rect 79 17 113 19
rect 79 -19 113 -17
rect 79 -104 113 -85
rect 175 85 209 104
rect 175 17 209 19
rect 175 -19 209 -17
rect 175 -104 209 -85
rect 271 85 305 104
rect 271 17 305 19
rect 271 -19 305 -17
rect 271 -104 305 -85
rect 367 85 401 104
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -104 401 -85
rect 463 85 497 104
rect 463 17 497 19
rect 463 -19 497 -17
rect 463 -104 497 -85
rect 577 85 611 119
rect 577 17 611 51
rect 577 -51 611 -17
rect 577 -119 611 -85
rect -611 -240 -577 -153
rect -465 -172 -449 -138
rect -415 -172 -399 -138
rect -273 -172 -257 -138
rect -223 -172 -207 -138
rect -81 -172 -65 -138
rect -31 -172 -15 -138
rect 111 -172 127 -138
rect 161 -172 177 -138
rect 303 -172 319 -138
rect 353 -172 369 -138
rect 577 -240 611 -153
rect -611 -274 -493 -240
rect -459 -274 -425 -240
rect -391 -274 -357 -240
rect -323 -274 -289 -240
rect -255 -274 -221 -240
rect -187 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 187 -240
rect 221 -274 255 -240
rect 289 -274 323 -240
rect 357 -274 391 -240
rect 425 -274 459 -240
rect 493 -274 611 -240
<< viali >>
rect -353 138 -319 172
rect -161 138 -127 172
rect 31 138 65 172
rect 223 138 257 172
rect 415 138 449 172
rect -497 51 -463 53
rect -497 19 -463 51
rect -497 -51 -463 -19
rect -497 -53 -463 -51
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -305 51 -271 53
rect -305 19 -271 51
rect -305 -51 -271 -19
rect -305 -53 -271 -51
rect -209 51 -175 53
rect -209 19 -175 51
rect -209 -51 -175 -19
rect -209 -53 -175 -51
rect -113 51 -79 53
rect -113 19 -79 51
rect -113 -51 -79 -19
rect -113 -53 -79 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 79 51 113 53
rect 79 19 113 51
rect 79 -51 113 -19
rect 79 -53 113 -51
rect 175 51 209 53
rect 175 19 209 51
rect 175 -51 209 -19
rect 175 -53 209 -51
rect 271 51 305 53
rect 271 19 305 51
rect 271 -51 305 -19
rect 271 -53 305 -51
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 463 51 497 53
rect 463 19 497 51
rect 463 -51 497 -19
rect 463 -53 497 -51
rect -449 -172 -415 -138
rect -257 -172 -223 -138
rect -65 -172 -31 -138
rect 127 -172 161 -138
rect 319 -172 353 -138
<< metal1 >>
rect -365 172 -307 178
rect -365 138 -353 172
rect -319 138 -307 172
rect -365 132 -307 138
rect -173 172 -115 178
rect -173 138 -161 172
rect -127 138 -115 172
rect -173 132 -115 138
rect 19 172 77 178
rect 19 138 31 172
rect 65 138 77 172
rect 19 132 77 138
rect 211 172 269 178
rect 211 138 223 172
rect 257 138 269 172
rect 211 132 269 138
rect 403 172 461 178
rect 403 138 415 172
rect 449 138 461 172
rect 403 132 461 138
rect -503 53 -457 100
rect -503 19 -497 53
rect -463 19 -457 53
rect -503 -19 -457 19
rect -503 -53 -497 -19
rect -463 -53 -457 -19
rect -503 -100 -457 -53
rect -407 53 -361 100
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -100 -361 -53
rect -311 53 -265 100
rect -311 19 -305 53
rect -271 19 -265 53
rect -311 -19 -265 19
rect -311 -53 -305 -19
rect -271 -53 -265 -19
rect -311 -100 -265 -53
rect -215 53 -169 100
rect -215 19 -209 53
rect -175 19 -169 53
rect -215 -19 -169 19
rect -215 -53 -209 -19
rect -175 -53 -169 -19
rect -215 -100 -169 -53
rect -119 53 -73 100
rect -119 19 -113 53
rect -79 19 -73 53
rect -119 -19 -73 19
rect -119 -53 -113 -19
rect -79 -53 -73 -19
rect -119 -100 -73 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 73 53 119 100
rect 73 19 79 53
rect 113 19 119 53
rect 73 -19 119 19
rect 73 -53 79 -19
rect 113 -53 119 -19
rect 73 -100 119 -53
rect 169 53 215 100
rect 169 19 175 53
rect 209 19 215 53
rect 169 -19 215 19
rect 169 -53 175 -19
rect 209 -53 215 -19
rect 169 -100 215 -53
rect 265 53 311 100
rect 265 19 271 53
rect 305 19 311 53
rect 265 -19 311 19
rect 265 -53 271 -19
rect 305 -53 311 -19
rect 265 -100 311 -53
rect 361 53 407 100
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -100 407 -53
rect 457 53 503 100
rect 457 19 463 53
rect 497 19 503 53
rect 457 -19 503 19
rect 457 -53 463 -19
rect 497 -53 503 -19
rect 457 -100 503 -53
rect -461 -138 -403 -132
rect -461 -172 -449 -138
rect -415 -172 -403 -138
rect -461 -178 -403 -172
rect -269 -138 -211 -132
rect -269 -172 -257 -138
rect -223 -172 -211 -138
rect -269 -178 -211 -172
rect -77 -138 -19 -132
rect -77 -172 -65 -138
rect -31 -172 -19 -138
rect -77 -178 -19 -172
rect 115 -138 173 -132
rect 115 -172 127 -138
rect 161 -172 173 -138
rect 115 -178 173 -172
rect 307 -138 365 -132
rect 307 -172 319 -138
rect 353 -172 365 -138
rect 307 -178 365 -172
<< properties >>
string FIXED_BBOX -594 -257 594 257
<< end >>
