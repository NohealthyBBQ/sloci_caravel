magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -1097 930 1097 1181
rect -1097 565 1097 816
rect -1097 200 1097 451
rect -1097 -165 1097 86
rect -1097 -530 1097 -279
rect -1097 -895 1097 -644
<< nwell >>
rect -1097 930 1097 1292
rect -1097 565 1097 927
rect -1097 200 1097 562
rect -1097 -165 1097 197
rect -1097 -530 1097 -168
rect -1097 -895 1097 -533
rect -1097 -1260 1097 -898
<< pmoslvt >>
rect -1003 1030 -803 1230
rect -745 1030 -545 1230
rect -487 1030 -287 1230
rect -229 1030 -29 1230
rect 29 1030 229 1230
rect 287 1030 487 1230
rect 545 1030 745 1230
rect 803 1030 1003 1230
rect -1003 665 -803 865
rect -745 665 -545 865
rect -487 665 -287 865
rect -229 665 -29 865
rect 29 665 229 865
rect 287 665 487 865
rect 545 665 745 865
rect 803 665 1003 865
rect -1003 300 -803 500
rect -745 300 -545 500
rect -487 300 -287 500
rect -229 300 -29 500
rect 29 300 229 500
rect 287 300 487 500
rect 545 300 745 500
rect 803 300 1003 500
rect -1003 -65 -803 135
rect -745 -65 -545 135
rect -487 -65 -287 135
rect -229 -65 -29 135
rect 29 -65 229 135
rect 287 -65 487 135
rect 545 -65 745 135
rect 803 -65 1003 135
rect -1003 -430 -803 -230
rect -745 -430 -545 -230
rect -487 -430 -287 -230
rect -229 -430 -29 -230
rect 29 -430 229 -230
rect 287 -430 487 -230
rect 545 -430 745 -230
rect 803 -430 1003 -230
rect -1003 -795 -803 -595
rect -745 -795 -545 -595
rect -487 -795 -287 -595
rect -229 -795 -29 -595
rect 29 -795 229 -595
rect 287 -795 487 -595
rect 545 -795 745 -595
rect 803 -795 1003 -595
rect -1003 -1160 -803 -960
rect -745 -1160 -545 -960
rect -487 -1160 -287 -960
rect -229 -1160 -29 -960
rect 29 -1160 229 -960
rect 287 -1160 487 -960
rect 545 -1160 745 -960
rect 803 -1160 1003 -960
<< pdiff >>
rect -1061 1215 -1003 1230
rect -1061 1181 -1049 1215
rect -1015 1181 -1003 1215
rect -1061 1147 -1003 1181
rect -1061 1113 -1049 1147
rect -1015 1113 -1003 1147
rect -1061 1079 -1003 1113
rect -1061 1045 -1049 1079
rect -1015 1045 -1003 1079
rect -1061 1030 -1003 1045
rect -803 1215 -745 1230
rect -803 1181 -791 1215
rect -757 1181 -745 1215
rect -803 1147 -745 1181
rect -803 1113 -791 1147
rect -757 1113 -745 1147
rect -803 1079 -745 1113
rect -803 1045 -791 1079
rect -757 1045 -745 1079
rect -803 1030 -745 1045
rect -545 1215 -487 1230
rect -545 1181 -533 1215
rect -499 1181 -487 1215
rect -545 1147 -487 1181
rect -545 1113 -533 1147
rect -499 1113 -487 1147
rect -545 1079 -487 1113
rect -545 1045 -533 1079
rect -499 1045 -487 1079
rect -545 1030 -487 1045
rect -287 1215 -229 1230
rect -287 1181 -275 1215
rect -241 1181 -229 1215
rect -287 1147 -229 1181
rect -287 1113 -275 1147
rect -241 1113 -229 1147
rect -287 1079 -229 1113
rect -287 1045 -275 1079
rect -241 1045 -229 1079
rect -287 1030 -229 1045
rect -29 1215 29 1230
rect -29 1181 -17 1215
rect 17 1181 29 1215
rect -29 1147 29 1181
rect -29 1113 -17 1147
rect 17 1113 29 1147
rect -29 1079 29 1113
rect -29 1045 -17 1079
rect 17 1045 29 1079
rect -29 1030 29 1045
rect 229 1215 287 1230
rect 229 1181 241 1215
rect 275 1181 287 1215
rect 229 1147 287 1181
rect 229 1113 241 1147
rect 275 1113 287 1147
rect 229 1079 287 1113
rect 229 1045 241 1079
rect 275 1045 287 1079
rect 229 1030 287 1045
rect 487 1215 545 1230
rect 487 1181 499 1215
rect 533 1181 545 1215
rect 487 1147 545 1181
rect 487 1113 499 1147
rect 533 1113 545 1147
rect 487 1079 545 1113
rect 487 1045 499 1079
rect 533 1045 545 1079
rect 487 1030 545 1045
rect 745 1215 803 1230
rect 745 1181 757 1215
rect 791 1181 803 1215
rect 745 1147 803 1181
rect 745 1113 757 1147
rect 791 1113 803 1147
rect 745 1079 803 1113
rect 745 1045 757 1079
rect 791 1045 803 1079
rect 745 1030 803 1045
rect 1003 1215 1061 1230
rect 1003 1181 1015 1215
rect 1049 1181 1061 1215
rect 1003 1147 1061 1181
rect 1003 1113 1015 1147
rect 1049 1113 1061 1147
rect 1003 1079 1061 1113
rect 1003 1045 1015 1079
rect 1049 1045 1061 1079
rect 1003 1030 1061 1045
rect -1061 850 -1003 865
rect -1061 816 -1049 850
rect -1015 816 -1003 850
rect -1061 782 -1003 816
rect -1061 748 -1049 782
rect -1015 748 -1003 782
rect -1061 714 -1003 748
rect -1061 680 -1049 714
rect -1015 680 -1003 714
rect -1061 665 -1003 680
rect -803 850 -745 865
rect -803 816 -791 850
rect -757 816 -745 850
rect -803 782 -745 816
rect -803 748 -791 782
rect -757 748 -745 782
rect -803 714 -745 748
rect -803 680 -791 714
rect -757 680 -745 714
rect -803 665 -745 680
rect -545 850 -487 865
rect -545 816 -533 850
rect -499 816 -487 850
rect -545 782 -487 816
rect -545 748 -533 782
rect -499 748 -487 782
rect -545 714 -487 748
rect -545 680 -533 714
rect -499 680 -487 714
rect -545 665 -487 680
rect -287 850 -229 865
rect -287 816 -275 850
rect -241 816 -229 850
rect -287 782 -229 816
rect -287 748 -275 782
rect -241 748 -229 782
rect -287 714 -229 748
rect -287 680 -275 714
rect -241 680 -229 714
rect -287 665 -229 680
rect -29 850 29 865
rect -29 816 -17 850
rect 17 816 29 850
rect -29 782 29 816
rect -29 748 -17 782
rect 17 748 29 782
rect -29 714 29 748
rect -29 680 -17 714
rect 17 680 29 714
rect -29 665 29 680
rect 229 850 287 865
rect 229 816 241 850
rect 275 816 287 850
rect 229 782 287 816
rect 229 748 241 782
rect 275 748 287 782
rect 229 714 287 748
rect 229 680 241 714
rect 275 680 287 714
rect 229 665 287 680
rect 487 850 545 865
rect 487 816 499 850
rect 533 816 545 850
rect 487 782 545 816
rect 487 748 499 782
rect 533 748 545 782
rect 487 714 545 748
rect 487 680 499 714
rect 533 680 545 714
rect 487 665 545 680
rect 745 850 803 865
rect 745 816 757 850
rect 791 816 803 850
rect 745 782 803 816
rect 745 748 757 782
rect 791 748 803 782
rect 745 714 803 748
rect 745 680 757 714
rect 791 680 803 714
rect 745 665 803 680
rect 1003 850 1061 865
rect 1003 816 1015 850
rect 1049 816 1061 850
rect 1003 782 1061 816
rect 1003 748 1015 782
rect 1049 748 1061 782
rect 1003 714 1061 748
rect 1003 680 1015 714
rect 1049 680 1061 714
rect 1003 665 1061 680
rect -1061 485 -1003 500
rect -1061 451 -1049 485
rect -1015 451 -1003 485
rect -1061 417 -1003 451
rect -1061 383 -1049 417
rect -1015 383 -1003 417
rect -1061 349 -1003 383
rect -1061 315 -1049 349
rect -1015 315 -1003 349
rect -1061 300 -1003 315
rect -803 485 -745 500
rect -803 451 -791 485
rect -757 451 -745 485
rect -803 417 -745 451
rect -803 383 -791 417
rect -757 383 -745 417
rect -803 349 -745 383
rect -803 315 -791 349
rect -757 315 -745 349
rect -803 300 -745 315
rect -545 485 -487 500
rect -545 451 -533 485
rect -499 451 -487 485
rect -545 417 -487 451
rect -545 383 -533 417
rect -499 383 -487 417
rect -545 349 -487 383
rect -545 315 -533 349
rect -499 315 -487 349
rect -545 300 -487 315
rect -287 485 -229 500
rect -287 451 -275 485
rect -241 451 -229 485
rect -287 417 -229 451
rect -287 383 -275 417
rect -241 383 -229 417
rect -287 349 -229 383
rect -287 315 -275 349
rect -241 315 -229 349
rect -287 300 -229 315
rect -29 485 29 500
rect -29 451 -17 485
rect 17 451 29 485
rect -29 417 29 451
rect -29 383 -17 417
rect 17 383 29 417
rect -29 349 29 383
rect -29 315 -17 349
rect 17 315 29 349
rect -29 300 29 315
rect 229 485 287 500
rect 229 451 241 485
rect 275 451 287 485
rect 229 417 287 451
rect 229 383 241 417
rect 275 383 287 417
rect 229 349 287 383
rect 229 315 241 349
rect 275 315 287 349
rect 229 300 287 315
rect 487 485 545 500
rect 487 451 499 485
rect 533 451 545 485
rect 487 417 545 451
rect 487 383 499 417
rect 533 383 545 417
rect 487 349 545 383
rect 487 315 499 349
rect 533 315 545 349
rect 487 300 545 315
rect 745 485 803 500
rect 745 451 757 485
rect 791 451 803 485
rect 745 417 803 451
rect 745 383 757 417
rect 791 383 803 417
rect 745 349 803 383
rect 745 315 757 349
rect 791 315 803 349
rect 745 300 803 315
rect 1003 485 1061 500
rect 1003 451 1015 485
rect 1049 451 1061 485
rect 1003 417 1061 451
rect 1003 383 1015 417
rect 1049 383 1061 417
rect 1003 349 1061 383
rect 1003 315 1015 349
rect 1049 315 1061 349
rect 1003 300 1061 315
rect -1061 120 -1003 135
rect -1061 86 -1049 120
rect -1015 86 -1003 120
rect -1061 52 -1003 86
rect -1061 18 -1049 52
rect -1015 18 -1003 52
rect -1061 -16 -1003 18
rect -1061 -50 -1049 -16
rect -1015 -50 -1003 -16
rect -1061 -65 -1003 -50
rect -803 120 -745 135
rect -803 86 -791 120
rect -757 86 -745 120
rect -803 52 -745 86
rect -803 18 -791 52
rect -757 18 -745 52
rect -803 -16 -745 18
rect -803 -50 -791 -16
rect -757 -50 -745 -16
rect -803 -65 -745 -50
rect -545 120 -487 135
rect -545 86 -533 120
rect -499 86 -487 120
rect -545 52 -487 86
rect -545 18 -533 52
rect -499 18 -487 52
rect -545 -16 -487 18
rect -545 -50 -533 -16
rect -499 -50 -487 -16
rect -545 -65 -487 -50
rect -287 120 -229 135
rect -287 86 -275 120
rect -241 86 -229 120
rect -287 52 -229 86
rect -287 18 -275 52
rect -241 18 -229 52
rect -287 -16 -229 18
rect -287 -50 -275 -16
rect -241 -50 -229 -16
rect -287 -65 -229 -50
rect -29 120 29 135
rect -29 86 -17 120
rect 17 86 29 120
rect -29 52 29 86
rect -29 18 -17 52
rect 17 18 29 52
rect -29 -16 29 18
rect -29 -50 -17 -16
rect 17 -50 29 -16
rect -29 -65 29 -50
rect 229 120 287 135
rect 229 86 241 120
rect 275 86 287 120
rect 229 52 287 86
rect 229 18 241 52
rect 275 18 287 52
rect 229 -16 287 18
rect 229 -50 241 -16
rect 275 -50 287 -16
rect 229 -65 287 -50
rect 487 120 545 135
rect 487 86 499 120
rect 533 86 545 120
rect 487 52 545 86
rect 487 18 499 52
rect 533 18 545 52
rect 487 -16 545 18
rect 487 -50 499 -16
rect 533 -50 545 -16
rect 487 -65 545 -50
rect 745 120 803 135
rect 745 86 757 120
rect 791 86 803 120
rect 745 52 803 86
rect 745 18 757 52
rect 791 18 803 52
rect 745 -16 803 18
rect 745 -50 757 -16
rect 791 -50 803 -16
rect 745 -65 803 -50
rect 1003 120 1061 135
rect 1003 86 1015 120
rect 1049 86 1061 120
rect 1003 52 1061 86
rect 1003 18 1015 52
rect 1049 18 1061 52
rect 1003 -16 1061 18
rect 1003 -50 1015 -16
rect 1049 -50 1061 -16
rect 1003 -65 1061 -50
rect -1061 -245 -1003 -230
rect -1061 -279 -1049 -245
rect -1015 -279 -1003 -245
rect -1061 -313 -1003 -279
rect -1061 -347 -1049 -313
rect -1015 -347 -1003 -313
rect -1061 -381 -1003 -347
rect -1061 -415 -1049 -381
rect -1015 -415 -1003 -381
rect -1061 -430 -1003 -415
rect -803 -245 -745 -230
rect -803 -279 -791 -245
rect -757 -279 -745 -245
rect -803 -313 -745 -279
rect -803 -347 -791 -313
rect -757 -347 -745 -313
rect -803 -381 -745 -347
rect -803 -415 -791 -381
rect -757 -415 -745 -381
rect -803 -430 -745 -415
rect -545 -245 -487 -230
rect -545 -279 -533 -245
rect -499 -279 -487 -245
rect -545 -313 -487 -279
rect -545 -347 -533 -313
rect -499 -347 -487 -313
rect -545 -381 -487 -347
rect -545 -415 -533 -381
rect -499 -415 -487 -381
rect -545 -430 -487 -415
rect -287 -245 -229 -230
rect -287 -279 -275 -245
rect -241 -279 -229 -245
rect -287 -313 -229 -279
rect -287 -347 -275 -313
rect -241 -347 -229 -313
rect -287 -381 -229 -347
rect -287 -415 -275 -381
rect -241 -415 -229 -381
rect -287 -430 -229 -415
rect -29 -245 29 -230
rect -29 -279 -17 -245
rect 17 -279 29 -245
rect -29 -313 29 -279
rect -29 -347 -17 -313
rect 17 -347 29 -313
rect -29 -381 29 -347
rect -29 -415 -17 -381
rect 17 -415 29 -381
rect -29 -430 29 -415
rect 229 -245 287 -230
rect 229 -279 241 -245
rect 275 -279 287 -245
rect 229 -313 287 -279
rect 229 -347 241 -313
rect 275 -347 287 -313
rect 229 -381 287 -347
rect 229 -415 241 -381
rect 275 -415 287 -381
rect 229 -430 287 -415
rect 487 -245 545 -230
rect 487 -279 499 -245
rect 533 -279 545 -245
rect 487 -313 545 -279
rect 487 -347 499 -313
rect 533 -347 545 -313
rect 487 -381 545 -347
rect 487 -415 499 -381
rect 533 -415 545 -381
rect 487 -430 545 -415
rect 745 -245 803 -230
rect 745 -279 757 -245
rect 791 -279 803 -245
rect 745 -313 803 -279
rect 745 -347 757 -313
rect 791 -347 803 -313
rect 745 -381 803 -347
rect 745 -415 757 -381
rect 791 -415 803 -381
rect 745 -430 803 -415
rect 1003 -245 1061 -230
rect 1003 -279 1015 -245
rect 1049 -279 1061 -245
rect 1003 -313 1061 -279
rect 1003 -347 1015 -313
rect 1049 -347 1061 -313
rect 1003 -381 1061 -347
rect 1003 -415 1015 -381
rect 1049 -415 1061 -381
rect 1003 -430 1061 -415
rect -1061 -610 -1003 -595
rect -1061 -644 -1049 -610
rect -1015 -644 -1003 -610
rect -1061 -678 -1003 -644
rect -1061 -712 -1049 -678
rect -1015 -712 -1003 -678
rect -1061 -746 -1003 -712
rect -1061 -780 -1049 -746
rect -1015 -780 -1003 -746
rect -1061 -795 -1003 -780
rect -803 -610 -745 -595
rect -803 -644 -791 -610
rect -757 -644 -745 -610
rect -803 -678 -745 -644
rect -803 -712 -791 -678
rect -757 -712 -745 -678
rect -803 -746 -745 -712
rect -803 -780 -791 -746
rect -757 -780 -745 -746
rect -803 -795 -745 -780
rect -545 -610 -487 -595
rect -545 -644 -533 -610
rect -499 -644 -487 -610
rect -545 -678 -487 -644
rect -545 -712 -533 -678
rect -499 -712 -487 -678
rect -545 -746 -487 -712
rect -545 -780 -533 -746
rect -499 -780 -487 -746
rect -545 -795 -487 -780
rect -287 -610 -229 -595
rect -287 -644 -275 -610
rect -241 -644 -229 -610
rect -287 -678 -229 -644
rect -287 -712 -275 -678
rect -241 -712 -229 -678
rect -287 -746 -229 -712
rect -287 -780 -275 -746
rect -241 -780 -229 -746
rect -287 -795 -229 -780
rect -29 -610 29 -595
rect -29 -644 -17 -610
rect 17 -644 29 -610
rect -29 -678 29 -644
rect -29 -712 -17 -678
rect 17 -712 29 -678
rect -29 -746 29 -712
rect -29 -780 -17 -746
rect 17 -780 29 -746
rect -29 -795 29 -780
rect 229 -610 287 -595
rect 229 -644 241 -610
rect 275 -644 287 -610
rect 229 -678 287 -644
rect 229 -712 241 -678
rect 275 -712 287 -678
rect 229 -746 287 -712
rect 229 -780 241 -746
rect 275 -780 287 -746
rect 229 -795 287 -780
rect 487 -610 545 -595
rect 487 -644 499 -610
rect 533 -644 545 -610
rect 487 -678 545 -644
rect 487 -712 499 -678
rect 533 -712 545 -678
rect 487 -746 545 -712
rect 487 -780 499 -746
rect 533 -780 545 -746
rect 487 -795 545 -780
rect 745 -610 803 -595
rect 745 -644 757 -610
rect 791 -644 803 -610
rect 745 -678 803 -644
rect 745 -712 757 -678
rect 791 -712 803 -678
rect 745 -746 803 -712
rect 745 -780 757 -746
rect 791 -780 803 -746
rect 745 -795 803 -780
rect 1003 -610 1061 -595
rect 1003 -644 1015 -610
rect 1049 -644 1061 -610
rect 1003 -678 1061 -644
rect 1003 -712 1015 -678
rect 1049 -712 1061 -678
rect 1003 -746 1061 -712
rect 1003 -780 1015 -746
rect 1049 -780 1061 -746
rect 1003 -795 1061 -780
rect -1061 -975 -1003 -960
rect -1061 -1009 -1049 -975
rect -1015 -1009 -1003 -975
rect -1061 -1043 -1003 -1009
rect -1061 -1077 -1049 -1043
rect -1015 -1077 -1003 -1043
rect -1061 -1111 -1003 -1077
rect -1061 -1145 -1049 -1111
rect -1015 -1145 -1003 -1111
rect -1061 -1160 -1003 -1145
rect -803 -975 -745 -960
rect -803 -1009 -791 -975
rect -757 -1009 -745 -975
rect -803 -1043 -745 -1009
rect -803 -1077 -791 -1043
rect -757 -1077 -745 -1043
rect -803 -1111 -745 -1077
rect -803 -1145 -791 -1111
rect -757 -1145 -745 -1111
rect -803 -1160 -745 -1145
rect -545 -975 -487 -960
rect -545 -1009 -533 -975
rect -499 -1009 -487 -975
rect -545 -1043 -487 -1009
rect -545 -1077 -533 -1043
rect -499 -1077 -487 -1043
rect -545 -1111 -487 -1077
rect -545 -1145 -533 -1111
rect -499 -1145 -487 -1111
rect -545 -1160 -487 -1145
rect -287 -975 -229 -960
rect -287 -1009 -275 -975
rect -241 -1009 -229 -975
rect -287 -1043 -229 -1009
rect -287 -1077 -275 -1043
rect -241 -1077 -229 -1043
rect -287 -1111 -229 -1077
rect -287 -1145 -275 -1111
rect -241 -1145 -229 -1111
rect -287 -1160 -229 -1145
rect -29 -975 29 -960
rect -29 -1009 -17 -975
rect 17 -1009 29 -975
rect -29 -1043 29 -1009
rect -29 -1077 -17 -1043
rect 17 -1077 29 -1043
rect -29 -1111 29 -1077
rect -29 -1145 -17 -1111
rect 17 -1145 29 -1111
rect -29 -1160 29 -1145
rect 229 -975 287 -960
rect 229 -1009 241 -975
rect 275 -1009 287 -975
rect 229 -1043 287 -1009
rect 229 -1077 241 -1043
rect 275 -1077 287 -1043
rect 229 -1111 287 -1077
rect 229 -1145 241 -1111
rect 275 -1145 287 -1111
rect 229 -1160 287 -1145
rect 487 -975 545 -960
rect 487 -1009 499 -975
rect 533 -1009 545 -975
rect 487 -1043 545 -1009
rect 487 -1077 499 -1043
rect 533 -1077 545 -1043
rect 487 -1111 545 -1077
rect 487 -1145 499 -1111
rect 533 -1145 545 -1111
rect 487 -1160 545 -1145
rect 745 -975 803 -960
rect 745 -1009 757 -975
rect 791 -1009 803 -975
rect 745 -1043 803 -1009
rect 745 -1077 757 -1043
rect 791 -1077 803 -1043
rect 745 -1111 803 -1077
rect 745 -1145 757 -1111
rect 791 -1145 803 -1111
rect 745 -1160 803 -1145
rect 1003 -975 1061 -960
rect 1003 -1009 1015 -975
rect 1049 -1009 1061 -975
rect 1003 -1043 1061 -1009
rect 1003 -1077 1015 -1043
rect 1049 -1077 1061 -1043
rect 1003 -1111 1061 -1077
rect 1003 -1145 1015 -1111
rect 1049 -1145 1061 -1111
rect 1003 -1160 1061 -1145
<< pdiffc >>
rect -1049 1181 -1015 1215
rect -1049 1113 -1015 1147
rect -1049 1045 -1015 1079
rect -791 1181 -757 1215
rect -791 1113 -757 1147
rect -791 1045 -757 1079
rect -533 1181 -499 1215
rect -533 1113 -499 1147
rect -533 1045 -499 1079
rect -275 1181 -241 1215
rect -275 1113 -241 1147
rect -275 1045 -241 1079
rect -17 1181 17 1215
rect -17 1113 17 1147
rect -17 1045 17 1079
rect 241 1181 275 1215
rect 241 1113 275 1147
rect 241 1045 275 1079
rect 499 1181 533 1215
rect 499 1113 533 1147
rect 499 1045 533 1079
rect 757 1181 791 1215
rect 757 1113 791 1147
rect 757 1045 791 1079
rect 1015 1181 1049 1215
rect 1015 1113 1049 1147
rect 1015 1045 1049 1079
rect -1049 816 -1015 850
rect -1049 748 -1015 782
rect -1049 680 -1015 714
rect -791 816 -757 850
rect -791 748 -757 782
rect -791 680 -757 714
rect -533 816 -499 850
rect -533 748 -499 782
rect -533 680 -499 714
rect -275 816 -241 850
rect -275 748 -241 782
rect -275 680 -241 714
rect -17 816 17 850
rect -17 748 17 782
rect -17 680 17 714
rect 241 816 275 850
rect 241 748 275 782
rect 241 680 275 714
rect 499 816 533 850
rect 499 748 533 782
rect 499 680 533 714
rect 757 816 791 850
rect 757 748 791 782
rect 757 680 791 714
rect 1015 816 1049 850
rect 1015 748 1049 782
rect 1015 680 1049 714
rect -1049 451 -1015 485
rect -1049 383 -1015 417
rect -1049 315 -1015 349
rect -791 451 -757 485
rect -791 383 -757 417
rect -791 315 -757 349
rect -533 451 -499 485
rect -533 383 -499 417
rect -533 315 -499 349
rect -275 451 -241 485
rect -275 383 -241 417
rect -275 315 -241 349
rect -17 451 17 485
rect -17 383 17 417
rect -17 315 17 349
rect 241 451 275 485
rect 241 383 275 417
rect 241 315 275 349
rect 499 451 533 485
rect 499 383 533 417
rect 499 315 533 349
rect 757 451 791 485
rect 757 383 791 417
rect 757 315 791 349
rect 1015 451 1049 485
rect 1015 383 1049 417
rect 1015 315 1049 349
rect -1049 86 -1015 120
rect -1049 18 -1015 52
rect -1049 -50 -1015 -16
rect -791 86 -757 120
rect -791 18 -757 52
rect -791 -50 -757 -16
rect -533 86 -499 120
rect -533 18 -499 52
rect -533 -50 -499 -16
rect -275 86 -241 120
rect -275 18 -241 52
rect -275 -50 -241 -16
rect -17 86 17 120
rect -17 18 17 52
rect -17 -50 17 -16
rect 241 86 275 120
rect 241 18 275 52
rect 241 -50 275 -16
rect 499 86 533 120
rect 499 18 533 52
rect 499 -50 533 -16
rect 757 86 791 120
rect 757 18 791 52
rect 757 -50 791 -16
rect 1015 86 1049 120
rect 1015 18 1049 52
rect 1015 -50 1049 -16
rect -1049 -279 -1015 -245
rect -1049 -347 -1015 -313
rect -1049 -415 -1015 -381
rect -791 -279 -757 -245
rect -791 -347 -757 -313
rect -791 -415 -757 -381
rect -533 -279 -499 -245
rect -533 -347 -499 -313
rect -533 -415 -499 -381
rect -275 -279 -241 -245
rect -275 -347 -241 -313
rect -275 -415 -241 -381
rect -17 -279 17 -245
rect -17 -347 17 -313
rect -17 -415 17 -381
rect 241 -279 275 -245
rect 241 -347 275 -313
rect 241 -415 275 -381
rect 499 -279 533 -245
rect 499 -347 533 -313
rect 499 -415 533 -381
rect 757 -279 791 -245
rect 757 -347 791 -313
rect 757 -415 791 -381
rect 1015 -279 1049 -245
rect 1015 -347 1049 -313
rect 1015 -415 1049 -381
rect -1049 -644 -1015 -610
rect -1049 -712 -1015 -678
rect -1049 -780 -1015 -746
rect -791 -644 -757 -610
rect -791 -712 -757 -678
rect -791 -780 -757 -746
rect -533 -644 -499 -610
rect -533 -712 -499 -678
rect -533 -780 -499 -746
rect -275 -644 -241 -610
rect -275 -712 -241 -678
rect -275 -780 -241 -746
rect -17 -644 17 -610
rect -17 -712 17 -678
rect -17 -780 17 -746
rect 241 -644 275 -610
rect 241 -712 275 -678
rect 241 -780 275 -746
rect 499 -644 533 -610
rect 499 -712 533 -678
rect 499 -780 533 -746
rect 757 -644 791 -610
rect 757 -712 791 -678
rect 757 -780 791 -746
rect 1015 -644 1049 -610
rect 1015 -712 1049 -678
rect 1015 -780 1049 -746
rect -1049 -1009 -1015 -975
rect -1049 -1077 -1015 -1043
rect -1049 -1145 -1015 -1111
rect -791 -1009 -757 -975
rect -791 -1077 -757 -1043
rect -791 -1145 -757 -1111
rect -533 -1009 -499 -975
rect -533 -1077 -499 -1043
rect -533 -1145 -499 -1111
rect -275 -1009 -241 -975
rect -275 -1077 -241 -1043
rect -275 -1145 -241 -1111
rect -17 -1009 17 -975
rect -17 -1077 17 -1043
rect -17 -1145 17 -1111
rect 241 -1009 275 -975
rect 241 -1077 275 -1043
rect 241 -1145 275 -1111
rect 499 -1009 533 -975
rect 499 -1077 533 -1043
rect 499 -1145 533 -1111
rect 757 -1009 791 -975
rect 757 -1077 791 -1043
rect 757 -1145 791 -1111
rect 1015 -1009 1049 -975
rect 1015 -1077 1049 -1043
rect 1015 -1145 1049 -1111
<< poly >>
rect -1003 1230 -803 1256
rect -745 1230 -545 1256
rect -487 1230 -287 1256
rect -229 1230 -29 1256
rect 29 1230 229 1256
rect 287 1230 487 1256
rect 545 1230 745 1256
rect 803 1230 1003 1256
rect -1003 983 -803 1030
rect -1003 949 -954 983
rect -920 949 -886 983
rect -852 949 -803 983
rect -1003 933 -803 949
rect -745 983 -545 1030
rect -745 949 -696 983
rect -662 949 -628 983
rect -594 949 -545 983
rect -745 933 -545 949
rect -487 983 -287 1030
rect -487 949 -438 983
rect -404 949 -370 983
rect -336 949 -287 983
rect -487 933 -287 949
rect -229 983 -29 1030
rect -229 949 -180 983
rect -146 949 -112 983
rect -78 949 -29 983
rect -229 933 -29 949
rect 29 983 229 1030
rect 29 949 78 983
rect 112 949 146 983
rect 180 949 229 983
rect 29 933 229 949
rect 287 983 487 1030
rect 287 949 336 983
rect 370 949 404 983
rect 438 949 487 983
rect 287 933 487 949
rect 545 983 745 1030
rect 545 949 594 983
rect 628 949 662 983
rect 696 949 745 983
rect 545 933 745 949
rect 803 983 1003 1030
rect 803 949 852 983
rect 886 949 920 983
rect 954 949 1003 983
rect 803 933 1003 949
rect -1003 865 -803 891
rect -745 865 -545 891
rect -487 865 -287 891
rect -229 865 -29 891
rect 29 865 229 891
rect 287 865 487 891
rect 545 865 745 891
rect 803 865 1003 891
rect -1003 618 -803 665
rect -1003 584 -954 618
rect -920 584 -886 618
rect -852 584 -803 618
rect -1003 568 -803 584
rect -745 618 -545 665
rect -745 584 -696 618
rect -662 584 -628 618
rect -594 584 -545 618
rect -745 568 -545 584
rect -487 618 -287 665
rect -487 584 -438 618
rect -404 584 -370 618
rect -336 584 -287 618
rect -487 568 -287 584
rect -229 618 -29 665
rect -229 584 -180 618
rect -146 584 -112 618
rect -78 584 -29 618
rect -229 568 -29 584
rect 29 618 229 665
rect 29 584 78 618
rect 112 584 146 618
rect 180 584 229 618
rect 29 568 229 584
rect 287 618 487 665
rect 287 584 336 618
rect 370 584 404 618
rect 438 584 487 618
rect 287 568 487 584
rect 545 618 745 665
rect 545 584 594 618
rect 628 584 662 618
rect 696 584 745 618
rect 545 568 745 584
rect 803 618 1003 665
rect 803 584 852 618
rect 886 584 920 618
rect 954 584 1003 618
rect 803 568 1003 584
rect -1003 500 -803 526
rect -745 500 -545 526
rect -487 500 -287 526
rect -229 500 -29 526
rect 29 500 229 526
rect 287 500 487 526
rect 545 500 745 526
rect 803 500 1003 526
rect -1003 253 -803 300
rect -1003 219 -954 253
rect -920 219 -886 253
rect -852 219 -803 253
rect -1003 203 -803 219
rect -745 253 -545 300
rect -745 219 -696 253
rect -662 219 -628 253
rect -594 219 -545 253
rect -745 203 -545 219
rect -487 253 -287 300
rect -487 219 -438 253
rect -404 219 -370 253
rect -336 219 -287 253
rect -487 203 -287 219
rect -229 253 -29 300
rect -229 219 -180 253
rect -146 219 -112 253
rect -78 219 -29 253
rect -229 203 -29 219
rect 29 253 229 300
rect 29 219 78 253
rect 112 219 146 253
rect 180 219 229 253
rect 29 203 229 219
rect 287 253 487 300
rect 287 219 336 253
rect 370 219 404 253
rect 438 219 487 253
rect 287 203 487 219
rect 545 253 745 300
rect 545 219 594 253
rect 628 219 662 253
rect 696 219 745 253
rect 545 203 745 219
rect 803 253 1003 300
rect 803 219 852 253
rect 886 219 920 253
rect 954 219 1003 253
rect 803 203 1003 219
rect -1003 135 -803 161
rect -745 135 -545 161
rect -487 135 -287 161
rect -229 135 -29 161
rect 29 135 229 161
rect 287 135 487 161
rect 545 135 745 161
rect 803 135 1003 161
rect -1003 -112 -803 -65
rect -1003 -146 -954 -112
rect -920 -146 -886 -112
rect -852 -146 -803 -112
rect -1003 -162 -803 -146
rect -745 -112 -545 -65
rect -745 -146 -696 -112
rect -662 -146 -628 -112
rect -594 -146 -545 -112
rect -745 -162 -545 -146
rect -487 -112 -287 -65
rect -487 -146 -438 -112
rect -404 -146 -370 -112
rect -336 -146 -287 -112
rect -487 -162 -287 -146
rect -229 -112 -29 -65
rect -229 -146 -180 -112
rect -146 -146 -112 -112
rect -78 -146 -29 -112
rect -229 -162 -29 -146
rect 29 -112 229 -65
rect 29 -146 78 -112
rect 112 -146 146 -112
rect 180 -146 229 -112
rect 29 -162 229 -146
rect 287 -112 487 -65
rect 287 -146 336 -112
rect 370 -146 404 -112
rect 438 -146 487 -112
rect 287 -162 487 -146
rect 545 -112 745 -65
rect 545 -146 594 -112
rect 628 -146 662 -112
rect 696 -146 745 -112
rect 545 -162 745 -146
rect 803 -112 1003 -65
rect 803 -146 852 -112
rect 886 -146 920 -112
rect 954 -146 1003 -112
rect 803 -162 1003 -146
rect -1003 -230 -803 -204
rect -745 -230 -545 -204
rect -487 -230 -287 -204
rect -229 -230 -29 -204
rect 29 -230 229 -204
rect 287 -230 487 -204
rect 545 -230 745 -204
rect 803 -230 1003 -204
rect -1003 -477 -803 -430
rect -1003 -511 -954 -477
rect -920 -511 -886 -477
rect -852 -511 -803 -477
rect -1003 -527 -803 -511
rect -745 -477 -545 -430
rect -745 -511 -696 -477
rect -662 -511 -628 -477
rect -594 -511 -545 -477
rect -745 -527 -545 -511
rect -487 -477 -287 -430
rect -487 -511 -438 -477
rect -404 -511 -370 -477
rect -336 -511 -287 -477
rect -487 -527 -287 -511
rect -229 -477 -29 -430
rect -229 -511 -180 -477
rect -146 -511 -112 -477
rect -78 -511 -29 -477
rect -229 -527 -29 -511
rect 29 -477 229 -430
rect 29 -511 78 -477
rect 112 -511 146 -477
rect 180 -511 229 -477
rect 29 -527 229 -511
rect 287 -477 487 -430
rect 287 -511 336 -477
rect 370 -511 404 -477
rect 438 -511 487 -477
rect 287 -527 487 -511
rect 545 -477 745 -430
rect 545 -511 594 -477
rect 628 -511 662 -477
rect 696 -511 745 -477
rect 545 -527 745 -511
rect 803 -477 1003 -430
rect 803 -511 852 -477
rect 886 -511 920 -477
rect 954 -511 1003 -477
rect 803 -527 1003 -511
rect -1003 -595 -803 -569
rect -745 -595 -545 -569
rect -487 -595 -287 -569
rect -229 -595 -29 -569
rect 29 -595 229 -569
rect 287 -595 487 -569
rect 545 -595 745 -569
rect 803 -595 1003 -569
rect -1003 -842 -803 -795
rect -1003 -876 -954 -842
rect -920 -876 -886 -842
rect -852 -876 -803 -842
rect -1003 -892 -803 -876
rect -745 -842 -545 -795
rect -745 -876 -696 -842
rect -662 -876 -628 -842
rect -594 -876 -545 -842
rect -745 -892 -545 -876
rect -487 -842 -287 -795
rect -487 -876 -438 -842
rect -404 -876 -370 -842
rect -336 -876 -287 -842
rect -487 -892 -287 -876
rect -229 -842 -29 -795
rect -229 -876 -180 -842
rect -146 -876 -112 -842
rect -78 -876 -29 -842
rect -229 -892 -29 -876
rect 29 -842 229 -795
rect 29 -876 78 -842
rect 112 -876 146 -842
rect 180 -876 229 -842
rect 29 -892 229 -876
rect 287 -842 487 -795
rect 287 -876 336 -842
rect 370 -876 404 -842
rect 438 -876 487 -842
rect 287 -892 487 -876
rect 545 -842 745 -795
rect 545 -876 594 -842
rect 628 -876 662 -842
rect 696 -876 745 -842
rect 545 -892 745 -876
rect 803 -842 1003 -795
rect 803 -876 852 -842
rect 886 -876 920 -842
rect 954 -876 1003 -842
rect 803 -892 1003 -876
rect -1003 -960 -803 -934
rect -745 -960 -545 -934
rect -487 -960 -287 -934
rect -229 -960 -29 -934
rect 29 -960 229 -934
rect 287 -960 487 -934
rect 545 -960 745 -934
rect 803 -960 1003 -934
rect -1003 -1207 -803 -1160
rect -1003 -1241 -954 -1207
rect -920 -1241 -886 -1207
rect -852 -1241 -803 -1207
rect -1003 -1257 -803 -1241
rect -745 -1207 -545 -1160
rect -745 -1241 -696 -1207
rect -662 -1241 -628 -1207
rect -594 -1241 -545 -1207
rect -745 -1257 -545 -1241
rect -487 -1207 -287 -1160
rect -487 -1241 -438 -1207
rect -404 -1241 -370 -1207
rect -336 -1241 -287 -1207
rect -487 -1257 -287 -1241
rect -229 -1207 -29 -1160
rect -229 -1241 -180 -1207
rect -146 -1241 -112 -1207
rect -78 -1241 -29 -1207
rect -229 -1257 -29 -1241
rect 29 -1207 229 -1160
rect 29 -1241 78 -1207
rect 112 -1241 146 -1207
rect 180 -1241 229 -1207
rect 29 -1257 229 -1241
rect 287 -1207 487 -1160
rect 287 -1241 336 -1207
rect 370 -1241 404 -1207
rect 438 -1241 487 -1207
rect 287 -1257 487 -1241
rect 545 -1207 745 -1160
rect 545 -1241 594 -1207
rect 628 -1241 662 -1207
rect 696 -1241 745 -1207
rect 545 -1257 745 -1241
rect 803 -1207 1003 -1160
rect 803 -1241 852 -1207
rect 886 -1241 920 -1207
rect 954 -1241 1003 -1207
rect 803 -1257 1003 -1241
<< polycont >>
rect -954 949 -920 983
rect -886 949 -852 983
rect -696 949 -662 983
rect -628 949 -594 983
rect -438 949 -404 983
rect -370 949 -336 983
rect -180 949 -146 983
rect -112 949 -78 983
rect 78 949 112 983
rect 146 949 180 983
rect 336 949 370 983
rect 404 949 438 983
rect 594 949 628 983
rect 662 949 696 983
rect 852 949 886 983
rect 920 949 954 983
rect -954 584 -920 618
rect -886 584 -852 618
rect -696 584 -662 618
rect -628 584 -594 618
rect -438 584 -404 618
rect -370 584 -336 618
rect -180 584 -146 618
rect -112 584 -78 618
rect 78 584 112 618
rect 146 584 180 618
rect 336 584 370 618
rect 404 584 438 618
rect 594 584 628 618
rect 662 584 696 618
rect 852 584 886 618
rect 920 584 954 618
rect -954 219 -920 253
rect -886 219 -852 253
rect -696 219 -662 253
rect -628 219 -594 253
rect -438 219 -404 253
rect -370 219 -336 253
rect -180 219 -146 253
rect -112 219 -78 253
rect 78 219 112 253
rect 146 219 180 253
rect 336 219 370 253
rect 404 219 438 253
rect 594 219 628 253
rect 662 219 696 253
rect 852 219 886 253
rect 920 219 954 253
rect -954 -146 -920 -112
rect -886 -146 -852 -112
rect -696 -146 -662 -112
rect -628 -146 -594 -112
rect -438 -146 -404 -112
rect -370 -146 -336 -112
rect -180 -146 -146 -112
rect -112 -146 -78 -112
rect 78 -146 112 -112
rect 146 -146 180 -112
rect 336 -146 370 -112
rect 404 -146 438 -112
rect 594 -146 628 -112
rect 662 -146 696 -112
rect 852 -146 886 -112
rect 920 -146 954 -112
rect -954 -511 -920 -477
rect -886 -511 -852 -477
rect -696 -511 -662 -477
rect -628 -511 -594 -477
rect -438 -511 -404 -477
rect -370 -511 -336 -477
rect -180 -511 -146 -477
rect -112 -511 -78 -477
rect 78 -511 112 -477
rect 146 -511 180 -477
rect 336 -511 370 -477
rect 404 -511 438 -477
rect 594 -511 628 -477
rect 662 -511 696 -477
rect 852 -511 886 -477
rect 920 -511 954 -477
rect -954 -876 -920 -842
rect -886 -876 -852 -842
rect -696 -876 -662 -842
rect -628 -876 -594 -842
rect -438 -876 -404 -842
rect -370 -876 -336 -842
rect -180 -876 -146 -842
rect -112 -876 -78 -842
rect 78 -876 112 -842
rect 146 -876 180 -842
rect 336 -876 370 -842
rect 404 -876 438 -842
rect 594 -876 628 -842
rect 662 -876 696 -842
rect 852 -876 886 -842
rect 920 -876 954 -842
rect -954 -1241 -920 -1207
rect -886 -1241 -852 -1207
rect -696 -1241 -662 -1207
rect -628 -1241 -594 -1207
rect -438 -1241 -404 -1207
rect -370 -1241 -336 -1207
rect -180 -1241 -146 -1207
rect -112 -1241 -78 -1207
rect 78 -1241 112 -1207
rect 146 -1241 180 -1207
rect 336 -1241 370 -1207
rect 404 -1241 438 -1207
rect 594 -1241 628 -1207
rect 662 -1241 696 -1207
rect 852 -1241 886 -1207
rect 920 -1241 954 -1207
<< locali >>
rect -1049 1215 -1015 1234
rect -1049 1147 -1015 1149
rect -1049 1111 -1015 1113
rect -1049 1026 -1015 1045
rect -791 1215 -757 1234
rect -791 1147 -757 1149
rect -791 1111 -757 1113
rect -791 1026 -757 1045
rect -533 1215 -499 1234
rect -533 1147 -499 1149
rect -533 1111 -499 1113
rect -533 1026 -499 1045
rect -275 1215 -241 1234
rect -275 1147 -241 1149
rect -275 1111 -241 1113
rect -275 1026 -241 1045
rect -17 1215 17 1234
rect -17 1147 17 1149
rect -17 1111 17 1113
rect -17 1026 17 1045
rect 241 1215 275 1234
rect 241 1147 275 1149
rect 241 1111 275 1113
rect 241 1026 275 1045
rect 499 1215 533 1234
rect 499 1147 533 1149
rect 499 1111 533 1113
rect 499 1026 533 1045
rect 757 1215 791 1234
rect 757 1147 791 1149
rect 757 1111 791 1113
rect 757 1026 791 1045
rect 1015 1215 1049 1234
rect 1015 1147 1049 1149
rect 1015 1111 1049 1113
rect 1015 1026 1049 1045
rect -1003 949 -956 983
rect -920 949 -886 983
rect -850 949 -803 983
rect -745 949 -698 983
rect -662 949 -628 983
rect -592 949 -545 983
rect -487 949 -440 983
rect -404 949 -370 983
rect -334 949 -287 983
rect -229 949 -182 983
rect -146 949 -112 983
rect -76 949 -29 983
rect 29 949 76 983
rect 112 949 146 983
rect 182 949 229 983
rect 287 949 334 983
rect 370 949 404 983
rect 440 949 487 983
rect 545 949 592 983
rect 628 949 662 983
rect 698 949 745 983
rect 803 949 850 983
rect 886 949 920 983
rect 956 949 1003 983
rect -1049 850 -1015 869
rect -1049 782 -1015 784
rect -1049 746 -1015 748
rect -1049 661 -1015 680
rect -791 850 -757 869
rect -791 782 -757 784
rect -791 746 -757 748
rect -791 661 -757 680
rect -533 850 -499 869
rect -533 782 -499 784
rect -533 746 -499 748
rect -533 661 -499 680
rect -275 850 -241 869
rect -275 782 -241 784
rect -275 746 -241 748
rect -275 661 -241 680
rect -17 850 17 869
rect -17 782 17 784
rect -17 746 17 748
rect -17 661 17 680
rect 241 850 275 869
rect 241 782 275 784
rect 241 746 275 748
rect 241 661 275 680
rect 499 850 533 869
rect 499 782 533 784
rect 499 746 533 748
rect 499 661 533 680
rect 757 850 791 869
rect 757 782 791 784
rect 757 746 791 748
rect 757 661 791 680
rect 1015 850 1049 869
rect 1015 782 1049 784
rect 1015 746 1049 748
rect 1015 661 1049 680
rect -1003 584 -956 618
rect -920 584 -886 618
rect -850 584 -803 618
rect -745 584 -698 618
rect -662 584 -628 618
rect -592 584 -545 618
rect -487 584 -440 618
rect -404 584 -370 618
rect -334 584 -287 618
rect -229 584 -182 618
rect -146 584 -112 618
rect -76 584 -29 618
rect 29 584 76 618
rect 112 584 146 618
rect 182 584 229 618
rect 287 584 334 618
rect 370 584 404 618
rect 440 584 487 618
rect 545 584 592 618
rect 628 584 662 618
rect 698 584 745 618
rect 803 584 850 618
rect 886 584 920 618
rect 956 584 1003 618
rect -1049 485 -1015 504
rect -1049 417 -1015 419
rect -1049 381 -1015 383
rect -1049 296 -1015 315
rect -791 485 -757 504
rect -791 417 -757 419
rect -791 381 -757 383
rect -791 296 -757 315
rect -533 485 -499 504
rect -533 417 -499 419
rect -533 381 -499 383
rect -533 296 -499 315
rect -275 485 -241 504
rect -275 417 -241 419
rect -275 381 -241 383
rect -275 296 -241 315
rect -17 485 17 504
rect -17 417 17 419
rect -17 381 17 383
rect -17 296 17 315
rect 241 485 275 504
rect 241 417 275 419
rect 241 381 275 383
rect 241 296 275 315
rect 499 485 533 504
rect 499 417 533 419
rect 499 381 533 383
rect 499 296 533 315
rect 757 485 791 504
rect 757 417 791 419
rect 757 381 791 383
rect 757 296 791 315
rect 1015 485 1049 504
rect 1015 417 1049 419
rect 1015 381 1049 383
rect 1015 296 1049 315
rect -1003 219 -956 253
rect -920 219 -886 253
rect -850 219 -803 253
rect -745 219 -698 253
rect -662 219 -628 253
rect -592 219 -545 253
rect -487 219 -440 253
rect -404 219 -370 253
rect -334 219 -287 253
rect -229 219 -182 253
rect -146 219 -112 253
rect -76 219 -29 253
rect 29 219 76 253
rect 112 219 146 253
rect 182 219 229 253
rect 287 219 334 253
rect 370 219 404 253
rect 440 219 487 253
rect 545 219 592 253
rect 628 219 662 253
rect 698 219 745 253
rect 803 219 850 253
rect 886 219 920 253
rect 956 219 1003 253
rect -1049 120 -1015 139
rect -1049 52 -1015 54
rect -1049 16 -1015 18
rect -1049 -69 -1015 -50
rect -791 120 -757 139
rect -791 52 -757 54
rect -791 16 -757 18
rect -791 -69 -757 -50
rect -533 120 -499 139
rect -533 52 -499 54
rect -533 16 -499 18
rect -533 -69 -499 -50
rect -275 120 -241 139
rect -275 52 -241 54
rect -275 16 -241 18
rect -275 -69 -241 -50
rect -17 120 17 139
rect -17 52 17 54
rect -17 16 17 18
rect -17 -69 17 -50
rect 241 120 275 139
rect 241 52 275 54
rect 241 16 275 18
rect 241 -69 275 -50
rect 499 120 533 139
rect 499 52 533 54
rect 499 16 533 18
rect 499 -69 533 -50
rect 757 120 791 139
rect 757 52 791 54
rect 757 16 791 18
rect 757 -69 791 -50
rect 1015 120 1049 139
rect 1015 52 1049 54
rect 1015 16 1049 18
rect 1015 -69 1049 -50
rect -1003 -146 -956 -112
rect -920 -146 -886 -112
rect -850 -146 -803 -112
rect -745 -146 -698 -112
rect -662 -146 -628 -112
rect -592 -146 -545 -112
rect -487 -146 -440 -112
rect -404 -146 -370 -112
rect -334 -146 -287 -112
rect -229 -146 -182 -112
rect -146 -146 -112 -112
rect -76 -146 -29 -112
rect 29 -146 76 -112
rect 112 -146 146 -112
rect 182 -146 229 -112
rect 287 -146 334 -112
rect 370 -146 404 -112
rect 440 -146 487 -112
rect 545 -146 592 -112
rect 628 -146 662 -112
rect 698 -146 745 -112
rect 803 -146 850 -112
rect 886 -146 920 -112
rect 956 -146 1003 -112
rect -1049 -245 -1015 -226
rect -1049 -313 -1015 -311
rect -1049 -349 -1015 -347
rect -1049 -434 -1015 -415
rect -791 -245 -757 -226
rect -791 -313 -757 -311
rect -791 -349 -757 -347
rect -791 -434 -757 -415
rect -533 -245 -499 -226
rect -533 -313 -499 -311
rect -533 -349 -499 -347
rect -533 -434 -499 -415
rect -275 -245 -241 -226
rect -275 -313 -241 -311
rect -275 -349 -241 -347
rect -275 -434 -241 -415
rect -17 -245 17 -226
rect -17 -313 17 -311
rect -17 -349 17 -347
rect -17 -434 17 -415
rect 241 -245 275 -226
rect 241 -313 275 -311
rect 241 -349 275 -347
rect 241 -434 275 -415
rect 499 -245 533 -226
rect 499 -313 533 -311
rect 499 -349 533 -347
rect 499 -434 533 -415
rect 757 -245 791 -226
rect 757 -313 791 -311
rect 757 -349 791 -347
rect 757 -434 791 -415
rect 1015 -245 1049 -226
rect 1015 -313 1049 -311
rect 1015 -349 1049 -347
rect 1015 -434 1049 -415
rect -1003 -511 -956 -477
rect -920 -511 -886 -477
rect -850 -511 -803 -477
rect -745 -511 -698 -477
rect -662 -511 -628 -477
rect -592 -511 -545 -477
rect -487 -511 -440 -477
rect -404 -511 -370 -477
rect -334 -511 -287 -477
rect -229 -511 -182 -477
rect -146 -511 -112 -477
rect -76 -511 -29 -477
rect 29 -511 76 -477
rect 112 -511 146 -477
rect 182 -511 229 -477
rect 287 -511 334 -477
rect 370 -511 404 -477
rect 440 -511 487 -477
rect 545 -511 592 -477
rect 628 -511 662 -477
rect 698 -511 745 -477
rect 803 -511 850 -477
rect 886 -511 920 -477
rect 956 -511 1003 -477
rect -1049 -610 -1015 -591
rect -1049 -678 -1015 -676
rect -1049 -714 -1015 -712
rect -1049 -799 -1015 -780
rect -791 -610 -757 -591
rect -791 -678 -757 -676
rect -791 -714 -757 -712
rect -791 -799 -757 -780
rect -533 -610 -499 -591
rect -533 -678 -499 -676
rect -533 -714 -499 -712
rect -533 -799 -499 -780
rect -275 -610 -241 -591
rect -275 -678 -241 -676
rect -275 -714 -241 -712
rect -275 -799 -241 -780
rect -17 -610 17 -591
rect -17 -678 17 -676
rect -17 -714 17 -712
rect -17 -799 17 -780
rect 241 -610 275 -591
rect 241 -678 275 -676
rect 241 -714 275 -712
rect 241 -799 275 -780
rect 499 -610 533 -591
rect 499 -678 533 -676
rect 499 -714 533 -712
rect 499 -799 533 -780
rect 757 -610 791 -591
rect 757 -678 791 -676
rect 757 -714 791 -712
rect 757 -799 791 -780
rect 1015 -610 1049 -591
rect 1015 -678 1049 -676
rect 1015 -714 1049 -712
rect 1015 -799 1049 -780
rect -1003 -876 -956 -842
rect -920 -876 -886 -842
rect -850 -876 -803 -842
rect -745 -876 -698 -842
rect -662 -876 -628 -842
rect -592 -876 -545 -842
rect -487 -876 -440 -842
rect -404 -876 -370 -842
rect -334 -876 -287 -842
rect -229 -876 -182 -842
rect -146 -876 -112 -842
rect -76 -876 -29 -842
rect 29 -876 76 -842
rect 112 -876 146 -842
rect 182 -876 229 -842
rect 287 -876 334 -842
rect 370 -876 404 -842
rect 440 -876 487 -842
rect 545 -876 592 -842
rect 628 -876 662 -842
rect 698 -876 745 -842
rect 803 -876 850 -842
rect 886 -876 920 -842
rect 956 -876 1003 -842
rect -1049 -975 -1015 -956
rect -1049 -1043 -1015 -1041
rect -1049 -1079 -1015 -1077
rect -1049 -1164 -1015 -1145
rect -791 -975 -757 -956
rect -791 -1043 -757 -1041
rect -791 -1079 -757 -1077
rect -791 -1164 -757 -1145
rect -533 -975 -499 -956
rect -533 -1043 -499 -1041
rect -533 -1079 -499 -1077
rect -533 -1164 -499 -1145
rect -275 -975 -241 -956
rect -275 -1043 -241 -1041
rect -275 -1079 -241 -1077
rect -275 -1164 -241 -1145
rect -17 -975 17 -956
rect -17 -1043 17 -1041
rect -17 -1079 17 -1077
rect -17 -1164 17 -1145
rect 241 -975 275 -956
rect 241 -1043 275 -1041
rect 241 -1079 275 -1077
rect 241 -1164 275 -1145
rect 499 -975 533 -956
rect 499 -1043 533 -1041
rect 499 -1079 533 -1077
rect 499 -1164 533 -1145
rect 757 -975 791 -956
rect 757 -1043 791 -1041
rect 757 -1079 791 -1077
rect 757 -1164 791 -1145
rect 1015 -975 1049 -956
rect 1015 -1043 1049 -1041
rect 1015 -1079 1049 -1077
rect 1015 -1164 1049 -1145
rect -1003 -1241 -956 -1207
rect -920 -1241 -886 -1207
rect -850 -1241 -803 -1207
rect -745 -1241 -698 -1207
rect -662 -1241 -628 -1207
rect -592 -1241 -545 -1207
rect -487 -1241 -440 -1207
rect -404 -1241 -370 -1207
rect -334 -1241 -287 -1207
rect -229 -1241 -182 -1207
rect -146 -1241 -112 -1207
rect -76 -1241 -29 -1207
rect 29 -1241 76 -1207
rect 112 -1241 146 -1207
rect 182 -1241 229 -1207
rect 287 -1241 334 -1207
rect 370 -1241 404 -1207
rect 440 -1241 487 -1207
rect 545 -1241 592 -1207
rect 628 -1241 662 -1207
rect 698 -1241 745 -1207
rect 803 -1241 850 -1207
rect 886 -1241 920 -1207
rect 956 -1241 1003 -1207
<< viali >>
rect -1049 1181 -1015 1183
rect -1049 1149 -1015 1181
rect -1049 1079 -1015 1111
rect -1049 1077 -1015 1079
rect -791 1181 -757 1183
rect -791 1149 -757 1181
rect -791 1079 -757 1111
rect -791 1077 -757 1079
rect -533 1181 -499 1183
rect -533 1149 -499 1181
rect -533 1079 -499 1111
rect -533 1077 -499 1079
rect -275 1181 -241 1183
rect -275 1149 -241 1181
rect -275 1079 -241 1111
rect -275 1077 -241 1079
rect -17 1181 17 1183
rect -17 1149 17 1181
rect -17 1079 17 1111
rect -17 1077 17 1079
rect 241 1181 275 1183
rect 241 1149 275 1181
rect 241 1079 275 1111
rect 241 1077 275 1079
rect 499 1181 533 1183
rect 499 1149 533 1181
rect 499 1079 533 1111
rect 499 1077 533 1079
rect 757 1181 791 1183
rect 757 1149 791 1181
rect 757 1079 791 1111
rect 757 1077 791 1079
rect 1015 1181 1049 1183
rect 1015 1149 1049 1181
rect 1015 1079 1049 1111
rect 1015 1077 1049 1079
rect -956 949 -954 983
rect -954 949 -922 983
rect -884 949 -852 983
rect -852 949 -850 983
rect -698 949 -696 983
rect -696 949 -664 983
rect -626 949 -594 983
rect -594 949 -592 983
rect -440 949 -438 983
rect -438 949 -406 983
rect -368 949 -336 983
rect -336 949 -334 983
rect -182 949 -180 983
rect -180 949 -148 983
rect -110 949 -78 983
rect -78 949 -76 983
rect 76 949 78 983
rect 78 949 110 983
rect 148 949 180 983
rect 180 949 182 983
rect 334 949 336 983
rect 336 949 368 983
rect 406 949 438 983
rect 438 949 440 983
rect 592 949 594 983
rect 594 949 626 983
rect 664 949 696 983
rect 696 949 698 983
rect 850 949 852 983
rect 852 949 884 983
rect 922 949 954 983
rect 954 949 956 983
rect -1049 816 -1015 818
rect -1049 784 -1015 816
rect -1049 714 -1015 746
rect -1049 712 -1015 714
rect -791 816 -757 818
rect -791 784 -757 816
rect -791 714 -757 746
rect -791 712 -757 714
rect -533 816 -499 818
rect -533 784 -499 816
rect -533 714 -499 746
rect -533 712 -499 714
rect -275 816 -241 818
rect -275 784 -241 816
rect -275 714 -241 746
rect -275 712 -241 714
rect -17 816 17 818
rect -17 784 17 816
rect -17 714 17 746
rect -17 712 17 714
rect 241 816 275 818
rect 241 784 275 816
rect 241 714 275 746
rect 241 712 275 714
rect 499 816 533 818
rect 499 784 533 816
rect 499 714 533 746
rect 499 712 533 714
rect 757 816 791 818
rect 757 784 791 816
rect 757 714 791 746
rect 757 712 791 714
rect 1015 816 1049 818
rect 1015 784 1049 816
rect 1015 714 1049 746
rect 1015 712 1049 714
rect -956 584 -954 618
rect -954 584 -922 618
rect -884 584 -852 618
rect -852 584 -850 618
rect -698 584 -696 618
rect -696 584 -664 618
rect -626 584 -594 618
rect -594 584 -592 618
rect -440 584 -438 618
rect -438 584 -406 618
rect -368 584 -336 618
rect -336 584 -334 618
rect -182 584 -180 618
rect -180 584 -148 618
rect -110 584 -78 618
rect -78 584 -76 618
rect 76 584 78 618
rect 78 584 110 618
rect 148 584 180 618
rect 180 584 182 618
rect 334 584 336 618
rect 336 584 368 618
rect 406 584 438 618
rect 438 584 440 618
rect 592 584 594 618
rect 594 584 626 618
rect 664 584 696 618
rect 696 584 698 618
rect 850 584 852 618
rect 852 584 884 618
rect 922 584 954 618
rect 954 584 956 618
rect -1049 451 -1015 453
rect -1049 419 -1015 451
rect -1049 349 -1015 381
rect -1049 347 -1015 349
rect -791 451 -757 453
rect -791 419 -757 451
rect -791 349 -757 381
rect -791 347 -757 349
rect -533 451 -499 453
rect -533 419 -499 451
rect -533 349 -499 381
rect -533 347 -499 349
rect -275 451 -241 453
rect -275 419 -241 451
rect -275 349 -241 381
rect -275 347 -241 349
rect -17 451 17 453
rect -17 419 17 451
rect -17 349 17 381
rect -17 347 17 349
rect 241 451 275 453
rect 241 419 275 451
rect 241 349 275 381
rect 241 347 275 349
rect 499 451 533 453
rect 499 419 533 451
rect 499 349 533 381
rect 499 347 533 349
rect 757 451 791 453
rect 757 419 791 451
rect 757 349 791 381
rect 757 347 791 349
rect 1015 451 1049 453
rect 1015 419 1049 451
rect 1015 349 1049 381
rect 1015 347 1049 349
rect -956 219 -954 253
rect -954 219 -922 253
rect -884 219 -852 253
rect -852 219 -850 253
rect -698 219 -696 253
rect -696 219 -664 253
rect -626 219 -594 253
rect -594 219 -592 253
rect -440 219 -438 253
rect -438 219 -406 253
rect -368 219 -336 253
rect -336 219 -334 253
rect -182 219 -180 253
rect -180 219 -148 253
rect -110 219 -78 253
rect -78 219 -76 253
rect 76 219 78 253
rect 78 219 110 253
rect 148 219 180 253
rect 180 219 182 253
rect 334 219 336 253
rect 336 219 368 253
rect 406 219 438 253
rect 438 219 440 253
rect 592 219 594 253
rect 594 219 626 253
rect 664 219 696 253
rect 696 219 698 253
rect 850 219 852 253
rect 852 219 884 253
rect 922 219 954 253
rect 954 219 956 253
rect -1049 86 -1015 88
rect -1049 54 -1015 86
rect -1049 -16 -1015 16
rect -1049 -18 -1015 -16
rect -791 86 -757 88
rect -791 54 -757 86
rect -791 -16 -757 16
rect -791 -18 -757 -16
rect -533 86 -499 88
rect -533 54 -499 86
rect -533 -16 -499 16
rect -533 -18 -499 -16
rect -275 86 -241 88
rect -275 54 -241 86
rect -275 -16 -241 16
rect -275 -18 -241 -16
rect -17 86 17 88
rect -17 54 17 86
rect -17 -16 17 16
rect -17 -18 17 -16
rect 241 86 275 88
rect 241 54 275 86
rect 241 -16 275 16
rect 241 -18 275 -16
rect 499 86 533 88
rect 499 54 533 86
rect 499 -16 533 16
rect 499 -18 533 -16
rect 757 86 791 88
rect 757 54 791 86
rect 757 -16 791 16
rect 757 -18 791 -16
rect 1015 86 1049 88
rect 1015 54 1049 86
rect 1015 -16 1049 16
rect 1015 -18 1049 -16
rect -956 -146 -954 -112
rect -954 -146 -922 -112
rect -884 -146 -852 -112
rect -852 -146 -850 -112
rect -698 -146 -696 -112
rect -696 -146 -664 -112
rect -626 -146 -594 -112
rect -594 -146 -592 -112
rect -440 -146 -438 -112
rect -438 -146 -406 -112
rect -368 -146 -336 -112
rect -336 -146 -334 -112
rect -182 -146 -180 -112
rect -180 -146 -148 -112
rect -110 -146 -78 -112
rect -78 -146 -76 -112
rect 76 -146 78 -112
rect 78 -146 110 -112
rect 148 -146 180 -112
rect 180 -146 182 -112
rect 334 -146 336 -112
rect 336 -146 368 -112
rect 406 -146 438 -112
rect 438 -146 440 -112
rect 592 -146 594 -112
rect 594 -146 626 -112
rect 664 -146 696 -112
rect 696 -146 698 -112
rect 850 -146 852 -112
rect 852 -146 884 -112
rect 922 -146 954 -112
rect 954 -146 956 -112
rect -1049 -279 -1015 -277
rect -1049 -311 -1015 -279
rect -1049 -381 -1015 -349
rect -1049 -383 -1015 -381
rect -791 -279 -757 -277
rect -791 -311 -757 -279
rect -791 -381 -757 -349
rect -791 -383 -757 -381
rect -533 -279 -499 -277
rect -533 -311 -499 -279
rect -533 -381 -499 -349
rect -533 -383 -499 -381
rect -275 -279 -241 -277
rect -275 -311 -241 -279
rect -275 -381 -241 -349
rect -275 -383 -241 -381
rect -17 -279 17 -277
rect -17 -311 17 -279
rect -17 -381 17 -349
rect -17 -383 17 -381
rect 241 -279 275 -277
rect 241 -311 275 -279
rect 241 -381 275 -349
rect 241 -383 275 -381
rect 499 -279 533 -277
rect 499 -311 533 -279
rect 499 -381 533 -349
rect 499 -383 533 -381
rect 757 -279 791 -277
rect 757 -311 791 -279
rect 757 -381 791 -349
rect 757 -383 791 -381
rect 1015 -279 1049 -277
rect 1015 -311 1049 -279
rect 1015 -381 1049 -349
rect 1015 -383 1049 -381
rect -956 -511 -954 -477
rect -954 -511 -922 -477
rect -884 -511 -852 -477
rect -852 -511 -850 -477
rect -698 -511 -696 -477
rect -696 -511 -664 -477
rect -626 -511 -594 -477
rect -594 -511 -592 -477
rect -440 -511 -438 -477
rect -438 -511 -406 -477
rect -368 -511 -336 -477
rect -336 -511 -334 -477
rect -182 -511 -180 -477
rect -180 -511 -148 -477
rect -110 -511 -78 -477
rect -78 -511 -76 -477
rect 76 -511 78 -477
rect 78 -511 110 -477
rect 148 -511 180 -477
rect 180 -511 182 -477
rect 334 -511 336 -477
rect 336 -511 368 -477
rect 406 -511 438 -477
rect 438 -511 440 -477
rect 592 -511 594 -477
rect 594 -511 626 -477
rect 664 -511 696 -477
rect 696 -511 698 -477
rect 850 -511 852 -477
rect 852 -511 884 -477
rect 922 -511 954 -477
rect 954 -511 956 -477
rect -1049 -644 -1015 -642
rect -1049 -676 -1015 -644
rect -1049 -746 -1015 -714
rect -1049 -748 -1015 -746
rect -791 -644 -757 -642
rect -791 -676 -757 -644
rect -791 -746 -757 -714
rect -791 -748 -757 -746
rect -533 -644 -499 -642
rect -533 -676 -499 -644
rect -533 -746 -499 -714
rect -533 -748 -499 -746
rect -275 -644 -241 -642
rect -275 -676 -241 -644
rect -275 -746 -241 -714
rect -275 -748 -241 -746
rect -17 -644 17 -642
rect -17 -676 17 -644
rect -17 -746 17 -714
rect -17 -748 17 -746
rect 241 -644 275 -642
rect 241 -676 275 -644
rect 241 -746 275 -714
rect 241 -748 275 -746
rect 499 -644 533 -642
rect 499 -676 533 -644
rect 499 -746 533 -714
rect 499 -748 533 -746
rect 757 -644 791 -642
rect 757 -676 791 -644
rect 757 -746 791 -714
rect 757 -748 791 -746
rect 1015 -644 1049 -642
rect 1015 -676 1049 -644
rect 1015 -746 1049 -714
rect 1015 -748 1049 -746
rect -956 -876 -954 -842
rect -954 -876 -922 -842
rect -884 -876 -852 -842
rect -852 -876 -850 -842
rect -698 -876 -696 -842
rect -696 -876 -664 -842
rect -626 -876 -594 -842
rect -594 -876 -592 -842
rect -440 -876 -438 -842
rect -438 -876 -406 -842
rect -368 -876 -336 -842
rect -336 -876 -334 -842
rect -182 -876 -180 -842
rect -180 -876 -148 -842
rect -110 -876 -78 -842
rect -78 -876 -76 -842
rect 76 -876 78 -842
rect 78 -876 110 -842
rect 148 -876 180 -842
rect 180 -876 182 -842
rect 334 -876 336 -842
rect 336 -876 368 -842
rect 406 -876 438 -842
rect 438 -876 440 -842
rect 592 -876 594 -842
rect 594 -876 626 -842
rect 664 -876 696 -842
rect 696 -876 698 -842
rect 850 -876 852 -842
rect 852 -876 884 -842
rect 922 -876 954 -842
rect 954 -876 956 -842
rect -1049 -1009 -1015 -1007
rect -1049 -1041 -1015 -1009
rect -1049 -1111 -1015 -1079
rect -1049 -1113 -1015 -1111
rect -791 -1009 -757 -1007
rect -791 -1041 -757 -1009
rect -791 -1111 -757 -1079
rect -791 -1113 -757 -1111
rect -533 -1009 -499 -1007
rect -533 -1041 -499 -1009
rect -533 -1111 -499 -1079
rect -533 -1113 -499 -1111
rect -275 -1009 -241 -1007
rect -275 -1041 -241 -1009
rect -275 -1111 -241 -1079
rect -275 -1113 -241 -1111
rect -17 -1009 17 -1007
rect -17 -1041 17 -1009
rect -17 -1111 17 -1079
rect -17 -1113 17 -1111
rect 241 -1009 275 -1007
rect 241 -1041 275 -1009
rect 241 -1111 275 -1079
rect 241 -1113 275 -1111
rect 499 -1009 533 -1007
rect 499 -1041 533 -1009
rect 499 -1111 533 -1079
rect 499 -1113 533 -1111
rect 757 -1009 791 -1007
rect 757 -1041 791 -1009
rect 757 -1111 791 -1079
rect 757 -1113 791 -1111
rect 1015 -1009 1049 -1007
rect 1015 -1041 1049 -1009
rect 1015 -1111 1049 -1079
rect 1015 -1113 1049 -1111
rect -956 -1241 -954 -1207
rect -954 -1241 -922 -1207
rect -884 -1241 -852 -1207
rect -852 -1241 -850 -1207
rect -698 -1241 -696 -1207
rect -696 -1241 -664 -1207
rect -626 -1241 -594 -1207
rect -594 -1241 -592 -1207
rect -440 -1241 -438 -1207
rect -438 -1241 -406 -1207
rect -368 -1241 -336 -1207
rect -336 -1241 -334 -1207
rect -182 -1241 -180 -1207
rect -180 -1241 -148 -1207
rect -110 -1241 -78 -1207
rect -78 -1241 -76 -1207
rect 76 -1241 78 -1207
rect 78 -1241 110 -1207
rect 148 -1241 180 -1207
rect 180 -1241 182 -1207
rect 334 -1241 336 -1207
rect 336 -1241 368 -1207
rect 406 -1241 438 -1207
rect 438 -1241 440 -1207
rect 592 -1241 594 -1207
rect 594 -1241 626 -1207
rect 664 -1241 696 -1207
rect 696 -1241 698 -1207
rect 850 -1241 852 -1207
rect 852 -1241 884 -1207
rect 922 -1241 954 -1207
rect 954 -1241 956 -1207
<< metal1 >>
rect -1055 1183 -1009 1230
rect -1055 1149 -1049 1183
rect -1015 1149 -1009 1183
rect -1055 1111 -1009 1149
rect -1055 1077 -1049 1111
rect -1015 1077 -1009 1111
rect -1055 1030 -1009 1077
rect -797 1183 -751 1230
rect -797 1149 -791 1183
rect -757 1149 -751 1183
rect -797 1111 -751 1149
rect -797 1077 -791 1111
rect -757 1077 -751 1111
rect -797 1030 -751 1077
rect -539 1183 -493 1230
rect -539 1149 -533 1183
rect -499 1149 -493 1183
rect -539 1111 -493 1149
rect -539 1077 -533 1111
rect -499 1077 -493 1111
rect -539 1030 -493 1077
rect -281 1183 -235 1230
rect -281 1149 -275 1183
rect -241 1149 -235 1183
rect -281 1111 -235 1149
rect -281 1077 -275 1111
rect -241 1077 -235 1111
rect -281 1030 -235 1077
rect -23 1183 23 1230
rect -23 1149 -17 1183
rect 17 1149 23 1183
rect -23 1111 23 1149
rect -23 1077 -17 1111
rect 17 1077 23 1111
rect -23 1030 23 1077
rect 235 1183 281 1230
rect 235 1149 241 1183
rect 275 1149 281 1183
rect 235 1111 281 1149
rect 235 1077 241 1111
rect 275 1077 281 1111
rect 235 1030 281 1077
rect 493 1183 539 1230
rect 493 1149 499 1183
rect 533 1149 539 1183
rect 493 1111 539 1149
rect 493 1077 499 1111
rect 533 1077 539 1111
rect 493 1030 539 1077
rect 751 1183 797 1230
rect 751 1149 757 1183
rect 791 1149 797 1183
rect 751 1111 797 1149
rect 751 1077 757 1111
rect 791 1077 797 1111
rect 751 1030 797 1077
rect 1009 1183 1055 1230
rect 1009 1149 1015 1183
rect 1049 1149 1055 1183
rect 1009 1111 1055 1149
rect 1009 1077 1015 1111
rect 1049 1077 1055 1111
rect 1009 1030 1055 1077
rect -999 983 -807 989
rect -999 949 -956 983
rect -922 949 -884 983
rect -850 949 -807 983
rect -999 943 -807 949
rect -741 983 -549 989
rect -741 949 -698 983
rect -664 949 -626 983
rect -592 949 -549 983
rect -741 943 -549 949
rect -483 983 -291 989
rect -483 949 -440 983
rect -406 949 -368 983
rect -334 949 -291 983
rect -483 943 -291 949
rect -225 983 -33 989
rect -225 949 -182 983
rect -148 949 -110 983
rect -76 949 -33 983
rect -225 943 -33 949
rect 33 983 225 989
rect 33 949 76 983
rect 110 949 148 983
rect 182 949 225 983
rect 33 943 225 949
rect 291 983 483 989
rect 291 949 334 983
rect 368 949 406 983
rect 440 949 483 983
rect 291 943 483 949
rect 549 983 741 989
rect 549 949 592 983
rect 626 949 664 983
rect 698 949 741 983
rect 549 943 741 949
rect 807 983 999 989
rect 807 949 850 983
rect 884 949 922 983
rect 956 949 999 983
rect 807 943 999 949
rect -1055 818 -1009 865
rect -1055 784 -1049 818
rect -1015 784 -1009 818
rect -1055 746 -1009 784
rect -1055 712 -1049 746
rect -1015 712 -1009 746
rect -1055 665 -1009 712
rect -797 818 -751 865
rect -797 784 -791 818
rect -757 784 -751 818
rect -797 746 -751 784
rect -797 712 -791 746
rect -757 712 -751 746
rect -797 665 -751 712
rect -539 818 -493 865
rect -539 784 -533 818
rect -499 784 -493 818
rect -539 746 -493 784
rect -539 712 -533 746
rect -499 712 -493 746
rect -539 665 -493 712
rect -281 818 -235 865
rect -281 784 -275 818
rect -241 784 -235 818
rect -281 746 -235 784
rect -281 712 -275 746
rect -241 712 -235 746
rect -281 665 -235 712
rect -23 818 23 865
rect -23 784 -17 818
rect 17 784 23 818
rect -23 746 23 784
rect -23 712 -17 746
rect 17 712 23 746
rect -23 665 23 712
rect 235 818 281 865
rect 235 784 241 818
rect 275 784 281 818
rect 235 746 281 784
rect 235 712 241 746
rect 275 712 281 746
rect 235 665 281 712
rect 493 818 539 865
rect 493 784 499 818
rect 533 784 539 818
rect 493 746 539 784
rect 493 712 499 746
rect 533 712 539 746
rect 493 665 539 712
rect 751 818 797 865
rect 751 784 757 818
rect 791 784 797 818
rect 751 746 797 784
rect 751 712 757 746
rect 791 712 797 746
rect 751 665 797 712
rect 1009 818 1055 865
rect 1009 784 1015 818
rect 1049 784 1055 818
rect 1009 746 1055 784
rect 1009 712 1015 746
rect 1049 712 1055 746
rect 1009 665 1055 712
rect -999 618 -807 624
rect -999 584 -956 618
rect -922 584 -884 618
rect -850 584 -807 618
rect -999 578 -807 584
rect -741 618 -549 624
rect -741 584 -698 618
rect -664 584 -626 618
rect -592 584 -549 618
rect -741 578 -549 584
rect -483 618 -291 624
rect -483 584 -440 618
rect -406 584 -368 618
rect -334 584 -291 618
rect -483 578 -291 584
rect -225 618 -33 624
rect -225 584 -182 618
rect -148 584 -110 618
rect -76 584 -33 618
rect -225 578 -33 584
rect 33 618 225 624
rect 33 584 76 618
rect 110 584 148 618
rect 182 584 225 618
rect 33 578 225 584
rect 291 618 483 624
rect 291 584 334 618
rect 368 584 406 618
rect 440 584 483 618
rect 291 578 483 584
rect 549 618 741 624
rect 549 584 592 618
rect 626 584 664 618
rect 698 584 741 618
rect 549 578 741 584
rect 807 618 999 624
rect 807 584 850 618
rect 884 584 922 618
rect 956 584 999 618
rect 807 578 999 584
rect -1055 453 -1009 500
rect -1055 419 -1049 453
rect -1015 419 -1009 453
rect -1055 381 -1009 419
rect -1055 347 -1049 381
rect -1015 347 -1009 381
rect -1055 300 -1009 347
rect -797 453 -751 500
rect -797 419 -791 453
rect -757 419 -751 453
rect -797 381 -751 419
rect -797 347 -791 381
rect -757 347 -751 381
rect -797 300 -751 347
rect -539 453 -493 500
rect -539 419 -533 453
rect -499 419 -493 453
rect -539 381 -493 419
rect -539 347 -533 381
rect -499 347 -493 381
rect -539 300 -493 347
rect -281 453 -235 500
rect -281 419 -275 453
rect -241 419 -235 453
rect -281 381 -235 419
rect -281 347 -275 381
rect -241 347 -235 381
rect -281 300 -235 347
rect -23 453 23 500
rect -23 419 -17 453
rect 17 419 23 453
rect -23 381 23 419
rect -23 347 -17 381
rect 17 347 23 381
rect -23 300 23 347
rect 235 453 281 500
rect 235 419 241 453
rect 275 419 281 453
rect 235 381 281 419
rect 235 347 241 381
rect 275 347 281 381
rect 235 300 281 347
rect 493 453 539 500
rect 493 419 499 453
rect 533 419 539 453
rect 493 381 539 419
rect 493 347 499 381
rect 533 347 539 381
rect 493 300 539 347
rect 751 453 797 500
rect 751 419 757 453
rect 791 419 797 453
rect 751 381 797 419
rect 751 347 757 381
rect 791 347 797 381
rect 751 300 797 347
rect 1009 453 1055 500
rect 1009 419 1015 453
rect 1049 419 1055 453
rect 1009 381 1055 419
rect 1009 347 1015 381
rect 1049 347 1055 381
rect 1009 300 1055 347
rect -999 253 -807 259
rect -999 219 -956 253
rect -922 219 -884 253
rect -850 219 -807 253
rect -999 213 -807 219
rect -741 253 -549 259
rect -741 219 -698 253
rect -664 219 -626 253
rect -592 219 -549 253
rect -741 213 -549 219
rect -483 253 -291 259
rect -483 219 -440 253
rect -406 219 -368 253
rect -334 219 -291 253
rect -483 213 -291 219
rect -225 253 -33 259
rect -225 219 -182 253
rect -148 219 -110 253
rect -76 219 -33 253
rect -225 213 -33 219
rect 33 253 225 259
rect 33 219 76 253
rect 110 219 148 253
rect 182 219 225 253
rect 33 213 225 219
rect 291 253 483 259
rect 291 219 334 253
rect 368 219 406 253
rect 440 219 483 253
rect 291 213 483 219
rect 549 253 741 259
rect 549 219 592 253
rect 626 219 664 253
rect 698 219 741 253
rect 549 213 741 219
rect 807 253 999 259
rect 807 219 850 253
rect 884 219 922 253
rect 956 219 999 253
rect 807 213 999 219
rect -1055 88 -1009 135
rect -1055 54 -1049 88
rect -1015 54 -1009 88
rect -1055 16 -1009 54
rect -1055 -18 -1049 16
rect -1015 -18 -1009 16
rect -1055 -65 -1009 -18
rect -797 88 -751 135
rect -797 54 -791 88
rect -757 54 -751 88
rect -797 16 -751 54
rect -797 -18 -791 16
rect -757 -18 -751 16
rect -797 -65 -751 -18
rect -539 88 -493 135
rect -539 54 -533 88
rect -499 54 -493 88
rect -539 16 -493 54
rect -539 -18 -533 16
rect -499 -18 -493 16
rect -539 -65 -493 -18
rect -281 88 -235 135
rect -281 54 -275 88
rect -241 54 -235 88
rect -281 16 -235 54
rect -281 -18 -275 16
rect -241 -18 -235 16
rect -281 -65 -235 -18
rect -23 88 23 135
rect -23 54 -17 88
rect 17 54 23 88
rect -23 16 23 54
rect -23 -18 -17 16
rect 17 -18 23 16
rect -23 -65 23 -18
rect 235 88 281 135
rect 235 54 241 88
rect 275 54 281 88
rect 235 16 281 54
rect 235 -18 241 16
rect 275 -18 281 16
rect 235 -65 281 -18
rect 493 88 539 135
rect 493 54 499 88
rect 533 54 539 88
rect 493 16 539 54
rect 493 -18 499 16
rect 533 -18 539 16
rect 493 -65 539 -18
rect 751 88 797 135
rect 751 54 757 88
rect 791 54 797 88
rect 751 16 797 54
rect 751 -18 757 16
rect 791 -18 797 16
rect 751 -65 797 -18
rect 1009 88 1055 135
rect 1009 54 1015 88
rect 1049 54 1055 88
rect 1009 16 1055 54
rect 1009 -18 1015 16
rect 1049 -18 1055 16
rect 1009 -65 1055 -18
rect -999 -112 -807 -106
rect -999 -146 -956 -112
rect -922 -146 -884 -112
rect -850 -146 -807 -112
rect -999 -152 -807 -146
rect -741 -112 -549 -106
rect -741 -146 -698 -112
rect -664 -146 -626 -112
rect -592 -146 -549 -112
rect -741 -152 -549 -146
rect -483 -112 -291 -106
rect -483 -146 -440 -112
rect -406 -146 -368 -112
rect -334 -146 -291 -112
rect -483 -152 -291 -146
rect -225 -112 -33 -106
rect -225 -146 -182 -112
rect -148 -146 -110 -112
rect -76 -146 -33 -112
rect -225 -152 -33 -146
rect 33 -112 225 -106
rect 33 -146 76 -112
rect 110 -146 148 -112
rect 182 -146 225 -112
rect 33 -152 225 -146
rect 291 -112 483 -106
rect 291 -146 334 -112
rect 368 -146 406 -112
rect 440 -146 483 -112
rect 291 -152 483 -146
rect 549 -112 741 -106
rect 549 -146 592 -112
rect 626 -146 664 -112
rect 698 -146 741 -112
rect 549 -152 741 -146
rect 807 -112 999 -106
rect 807 -146 850 -112
rect 884 -146 922 -112
rect 956 -146 999 -112
rect 807 -152 999 -146
rect -1055 -277 -1009 -230
rect -1055 -311 -1049 -277
rect -1015 -311 -1009 -277
rect -1055 -349 -1009 -311
rect -1055 -383 -1049 -349
rect -1015 -383 -1009 -349
rect -1055 -430 -1009 -383
rect -797 -277 -751 -230
rect -797 -311 -791 -277
rect -757 -311 -751 -277
rect -797 -349 -751 -311
rect -797 -383 -791 -349
rect -757 -383 -751 -349
rect -797 -430 -751 -383
rect -539 -277 -493 -230
rect -539 -311 -533 -277
rect -499 -311 -493 -277
rect -539 -349 -493 -311
rect -539 -383 -533 -349
rect -499 -383 -493 -349
rect -539 -430 -493 -383
rect -281 -277 -235 -230
rect -281 -311 -275 -277
rect -241 -311 -235 -277
rect -281 -349 -235 -311
rect -281 -383 -275 -349
rect -241 -383 -235 -349
rect -281 -430 -235 -383
rect -23 -277 23 -230
rect -23 -311 -17 -277
rect 17 -311 23 -277
rect -23 -349 23 -311
rect -23 -383 -17 -349
rect 17 -383 23 -349
rect -23 -430 23 -383
rect 235 -277 281 -230
rect 235 -311 241 -277
rect 275 -311 281 -277
rect 235 -349 281 -311
rect 235 -383 241 -349
rect 275 -383 281 -349
rect 235 -430 281 -383
rect 493 -277 539 -230
rect 493 -311 499 -277
rect 533 -311 539 -277
rect 493 -349 539 -311
rect 493 -383 499 -349
rect 533 -383 539 -349
rect 493 -430 539 -383
rect 751 -277 797 -230
rect 751 -311 757 -277
rect 791 -311 797 -277
rect 751 -349 797 -311
rect 751 -383 757 -349
rect 791 -383 797 -349
rect 751 -430 797 -383
rect 1009 -277 1055 -230
rect 1009 -311 1015 -277
rect 1049 -311 1055 -277
rect 1009 -349 1055 -311
rect 1009 -383 1015 -349
rect 1049 -383 1055 -349
rect 1009 -430 1055 -383
rect -999 -477 -807 -471
rect -999 -511 -956 -477
rect -922 -511 -884 -477
rect -850 -511 -807 -477
rect -999 -517 -807 -511
rect -741 -477 -549 -471
rect -741 -511 -698 -477
rect -664 -511 -626 -477
rect -592 -511 -549 -477
rect -741 -517 -549 -511
rect -483 -477 -291 -471
rect -483 -511 -440 -477
rect -406 -511 -368 -477
rect -334 -511 -291 -477
rect -483 -517 -291 -511
rect -225 -477 -33 -471
rect -225 -511 -182 -477
rect -148 -511 -110 -477
rect -76 -511 -33 -477
rect -225 -517 -33 -511
rect 33 -477 225 -471
rect 33 -511 76 -477
rect 110 -511 148 -477
rect 182 -511 225 -477
rect 33 -517 225 -511
rect 291 -477 483 -471
rect 291 -511 334 -477
rect 368 -511 406 -477
rect 440 -511 483 -477
rect 291 -517 483 -511
rect 549 -477 741 -471
rect 549 -511 592 -477
rect 626 -511 664 -477
rect 698 -511 741 -477
rect 549 -517 741 -511
rect 807 -477 999 -471
rect 807 -511 850 -477
rect 884 -511 922 -477
rect 956 -511 999 -477
rect 807 -517 999 -511
rect -1055 -642 -1009 -595
rect -1055 -676 -1049 -642
rect -1015 -676 -1009 -642
rect -1055 -714 -1009 -676
rect -1055 -748 -1049 -714
rect -1015 -748 -1009 -714
rect -1055 -795 -1009 -748
rect -797 -642 -751 -595
rect -797 -676 -791 -642
rect -757 -676 -751 -642
rect -797 -714 -751 -676
rect -797 -748 -791 -714
rect -757 -748 -751 -714
rect -797 -795 -751 -748
rect -539 -642 -493 -595
rect -539 -676 -533 -642
rect -499 -676 -493 -642
rect -539 -714 -493 -676
rect -539 -748 -533 -714
rect -499 -748 -493 -714
rect -539 -795 -493 -748
rect -281 -642 -235 -595
rect -281 -676 -275 -642
rect -241 -676 -235 -642
rect -281 -714 -235 -676
rect -281 -748 -275 -714
rect -241 -748 -235 -714
rect -281 -795 -235 -748
rect -23 -642 23 -595
rect -23 -676 -17 -642
rect 17 -676 23 -642
rect -23 -714 23 -676
rect -23 -748 -17 -714
rect 17 -748 23 -714
rect -23 -795 23 -748
rect 235 -642 281 -595
rect 235 -676 241 -642
rect 275 -676 281 -642
rect 235 -714 281 -676
rect 235 -748 241 -714
rect 275 -748 281 -714
rect 235 -795 281 -748
rect 493 -642 539 -595
rect 493 -676 499 -642
rect 533 -676 539 -642
rect 493 -714 539 -676
rect 493 -748 499 -714
rect 533 -748 539 -714
rect 493 -795 539 -748
rect 751 -642 797 -595
rect 751 -676 757 -642
rect 791 -676 797 -642
rect 751 -714 797 -676
rect 751 -748 757 -714
rect 791 -748 797 -714
rect 751 -795 797 -748
rect 1009 -642 1055 -595
rect 1009 -676 1015 -642
rect 1049 -676 1055 -642
rect 1009 -714 1055 -676
rect 1009 -748 1015 -714
rect 1049 -748 1055 -714
rect 1009 -795 1055 -748
rect -999 -842 -807 -836
rect -999 -876 -956 -842
rect -922 -876 -884 -842
rect -850 -876 -807 -842
rect -999 -882 -807 -876
rect -741 -842 -549 -836
rect -741 -876 -698 -842
rect -664 -876 -626 -842
rect -592 -876 -549 -842
rect -741 -882 -549 -876
rect -483 -842 -291 -836
rect -483 -876 -440 -842
rect -406 -876 -368 -842
rect -334 -876 -291 -842
rect -483 -882 -291 -876
rect -225 -842 -33 -836
rect -225 -876 -182 -842
rect -148 -876 -110 -842
rect -76 -876 -33 -842
rect -225 -882 -33 -876
rect 33 -842 225 -836
rect 33 -876 76 -842
rect 110 -876 148 -842
rect 182 -876 225 -842
rect 33 -882 225 -876
rect 291 -842 483 -836
rect 291 -876 334 -842
rect 368 -876 406 -842
rect 440 -876 483 -842
rect 291 -882 483 -876
rect 549 -842 741 -836
rect 549 -876 592 -842
rect 626 -876 664 -842
rect 698 -876 741 -842
rect 549 -882 741 -876
rect 807 -842 999 -836
rect 807 -876 850 -842
rect 884 -876 922 -842
rect 956 -876 999 -842
rect 807 -882 999 -876
rect -1055 -1007 -1009 -960
rect -1055 -1041 -1049 -1007
rect -1015 -1041 -1009 -1007
rect -1055 -1079 -1009 -1041
rect -1055 -1113 -1049 -1079
rect -1015 -1113 -1009 -1079
rect -1055 -1160 -1009 -1113
rect -797 -1007 -751 -960
rect -797 -1041 -791 -1007
rect -757 -1041 -751 -1007
rect -797 -1079 -751 -1041
rect -797 -1113 -791 -1079
rect -757 -1113 -751 -1079
rect -797 -1160 -751 -1113
rect -539 -1007 -493 -960
rect -539 -1041 -533 -1007
rect -499 -1041 -493 -1007
rect -539 -1079 -493 -1041
rect -539 -1113 -533 -1079
rect -499 -1113 -493 -1079
rect -539 -1160 -493 -1113
rect -281 -1007 -235 -960
rect -281 -1041 -275 -1007
rect -241 -1041 -235 -1007
rect -281 -1079 -235 -1041
rect -281 -1113 -275 -1079
rect -241 -1113 -235 -1079
rect -281 -1160 -235 -1113
rect -23 -1007 23 -960
rect -23 -1041 -17 -1007
rect 17 -1041 23 -1007
rect -23 -1079 23 -1041
rect -23 -1113 -17 -1079
rect 17 -1113 23 -1079
rect -23 -1160 23 -1113
rect 235 -1007 281 -960
rect 235 -1041 241 -1007
rect 275 -1041 281 -1007
rect 235 -1079 281 -1041
rect 235 -1113 241 -1079
rect 275 -1113 281 -1079
rect 235 -1160 281 -1113
rect 493 -1007 539 -960
rect 493 -1041 499 -1007
rect 533 -1041 539 -1007
rect 493 -1079 539 -1041
rect 493 -1113 499 -1079
rect 533 -1113 539 -1079
rect 493 -1160 539 -1113
rect 751 -1007 797 -960
rect 751 -1041 757 -1007
rect 791 -1041 797 -1007
rect 751 -1079 797 -1041
rect 751 -1113 757 -1079
rect 791 -1113 797 -1079
rect 751 -1160 797 -1113
rect 1009 -1007 1055 -960
rect 1009 -1041 1015 -1007
rect 1049 -1041 1055 -1007
rect 1009 -1079 1055 -1041
rect 1009 -1113 1015 -1079
rect 1049 -1113 1055 -1079
rect 1009 -1160 1055 -1113
rect -999 -1207 -807 -1201
rect -999 -1241 -956 -1207
rect -922 -1241 -884 -1207
rect -850 -1241 -807 -1207
rect -999 -1247 -807 -1241
rect -741 -1207 -549 -1201
rect -741 -1241 -698 -1207
rect -664 -1241 -626 -1207
rect -592 -1241 -549 -1207
rect -741 -1247 -549 -1241
rect -483 -1207 -291 -1201
rect -483 -1241 -440 -1207
rect -406 -1241 -368 -1207
rect -334 -1241 -291 -1207
rect -483 -1247 -291 -1241
rect -225 -1207 -33 -1201
rect -225 -1241 -182 -1207
rect -148 -1241 -110 -1207
rect -76 -1241 -33 -1207
rect -225 -1247 -33 -1241
rect 33 -1207 225 -1201
rect 33 -1241 76 -1207
rect 110 -1241 148 -1207
rect 182 -1241 225 -1207
rect 33 -1247 225 -1241
rect 291 -1207 483 -1201
rect 291 -1241 334 -1207
rect 368 -1241 406 -1207
rect 440 -1241 483 -1207
rect 291 -1247 483 -1241
rect 549 -1207 741 -1201
rect 549 -1241 592 -1207
rect 626 -1241 664 -1207
rect 698 -1241 741 -1207
rect 549 -1247 741 -1241
rect 807 -1207 999 -1201
rect 807 -1241 850 -1207
rect 884 -1241 922 -1207
rect 956 -1241 999 -1207
rect 807 -1247 999 -1241
<< end >>
