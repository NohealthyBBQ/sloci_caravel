magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 4525 -40 4560 105
rect 5040 -40 5075 105
rect 4525 -660 4560 -515
rect 5040 -655 5075 -510
rect 4525 -1155 4560 -1045
rect 4250 -1190 4560 -1155
rect 5040 -1185 5075 -1040
rect 4250 -1303 4560 -1285
rect 4250 -1337 4352 -1303
rect 4386 -1337 4424 -1303
rect 4458 -1337 4560 -1303
rect 4250 -1355 4560 -1337
rect 4250 -1505 4560 -1470
<< viali >>
rect 4352 -1337 4386 -1303
rect 4424 -1337 4458 -1303
<< metal1 >>
rect 3300 860 5110 920
rect 4610 300 4670 860
rect 4700 806 4780 820
rect 4700 754 4714 806
rect 4766 800 4780 806
rect 4766 754 4900 800
rect 4700 750 4900 754
rect 4700 740 4780 750
rect 4820 706 4900 720
rect 4820 700 4834 706
rect 4700 654 4834 700
rect 4886 654 4900 706
rect 4700 650 4900 654
rect 4820 640 4900 650
rect 4700 606 4780 620
rect 4700 554 4714 606
rect 4766 600 4780 606
rect 4766 560 4900 600
rect 4766 554 4780 560
rect 4700 540 4780 554
rect 4820 510 4900 520
rect 4700 506 4900 510
rect 4700 460 4834 506
rect 4820 454 4834 460
rect 4886 454 4900 506
rect 4820 440 4900 454
rect 4700 416 4780 430
rect 4700 364 4714 416
rect 4766 410 4780 416
rect 4766 370 4900 410
rect 4766 364 4780 370
rect 4700 350 4780 364
rect 4820 320 4900 330
rect 4700 316 4900 320
rect 4700 270 4834 316
rect 4820 264 4834 270
rect 4886 264 4900 316
rect 4820 250 4900 264
rect 4700 220 4780 230
rect 4700 216 4900 220
rect 4700 164 4714 216
rect 4766 170 4900 216
rect 4930 210 4990 860
rect 4766 164 4780 170
rect 4700 150 4780 164
rect 3300 -50 5110 10
rect 4610 -410 4670 -50
rect 4700 -114 4780 -100
rect 4700 -166 4714 -114
rect 4766 -166 4780 -114
rect 4700 -180 4780 -166
rect 4820 -204 4900 -190
rect 4820 -256 4834 -204
rect 4886 -256 4900 -204
rect 4820 -270 4900 -256
rect 4700 -304 4780 -290
rect 4700 -356 4714 -304
rect 4766 -356 4780 -304
rect 4930 -310 4990 -50
rect 4700 -370 4780 -356
rect 4820 -394 4900 -380
rect 4820 -446 4834 -394
rect 4886 -446 4900 -394
rect 4820 -460 4900 -446
rect 3300 -640 5110 -580
rect 4610 -670 4990 -640
rect 4610 -830 4670 -670
rect 4700 -724 4780 -710
rect 4700 -776 4714 -724
rect 4766 -776 4780 -724
rect 4700 -790 4780 -776
rect 4820 -824 4900 -810
rect 4820 -876 4834 -824
rect 4886 -876 4900 -824
rect 4820 -890 4900 -876
rect 4700 -914 4780 -900
rect 4700 -966 4714 -914
rect 4766 -966 4780 -914
rect 4930 -930 4990 -670
rect 4700 -980 4780 -966
rect 3300 -1180 5110 -1120
rect 3910 -1254 3990 -1240
rect 3820 -1360 3880 -1290
rect 3910 -1306 3924 -1254
rect 3976 -1262 3990 -1254
rect 4700 -1254 4780 -1240
rect 3976 -1306 4110 -1262
rect 3910 -1308 4110 -1306
rect 3910 -1320 3990 -1308
rect 4030 -1350 4110 -1340
rect 3910 -1354 4110 -1350
rect 3910 -1396 4044 -1354
rect 4030 -1406 4044 -1396
rect 4096 -1406 4110 -1354
rect 4030 -1420 4110 -1406
rect 4140 -1480 4200 -1290
rect 4320 -1294 4490 -1285
rect 4320 -1346 4347 -1294
rect 4399 -1346 4411 -1294
rect 4463 -1346 4490 -1294
rect 4320 -1355 4490 -1346
rect 4610 -1360 4670 -1290
rect 4700 -1306 4714 -1254
rect 4766 -1306 4780 -1254
rect 4700 -1320 4780 -1306
rect 4820 -1354 4900 -1340
rect 4820 -1406 4834 -1354
rect 4886 -1406 4900 -1354
rect 4930 -1360 4990 -1180
rect 4820 -1420 4900 -1406
rect 3300 -1540 5110 -1480
<< via1 >>
rect 4714 754 4766 806
rect 4834 654 4886 706
rect 4714 554 4766 606
rect 4834 454 4886 506
rect 4714 364 4766 416
rect 4834 264 4886 316
rect 4714 164 4766 216
rect 4714 -166 4766 -114
rect 4834 -256 4886 -204
rect 4714 -356 4766 -304
rect 4834 -446 4886 -394
rect 4714 -776 4766 -724
rect 4834 -876 4886 -824
rect 4714 -966 4766 -914
rect 3924 -1306 3976 -1254
rect 4044 -1406 4096 -1354
rect 4347 -1303 4399 -1294
rect 4347 -1337 4352 -1303
rect 4352 -1337 4386 -1303
rect 4386 -1337 4399 -1303
rect 4347 -1346 4399 -1337
rect 4411 -1303 4463 -1294
rect 4411 -1337 4424 -1303
rect 4424 -1337 4458 -1303
rect 4458 -1337 4463 -1303
rect 4411 -1346 4463 -1337
rect 4714 -1306 4766 -1254
rect 4834 -1406 4886 -1354
<< metal2 >>
rect 4520 806 4780 920
rect 4950 910 5110 920
rect 4520 754 4714 806
rect 4766 754 4780 806
rect 4520 606 4780 754
rect 4520 554 4714 606
rect 4766 554 4780 606
rect 4520 416 4780 554
rect 4520 364 4714 416
rect 4766 364 4780 416
rect 4520 216 4780 364
rect 4520 164 4714 216
rect 4766 164 4780 216
rect 4520 -114 4780 164
rect 4820 888 5110 910
rect 4820 832 5002 888
rect 5058 832 5110 888
rect 4820 808 5110 832
rect 4820 752 5002 808
rect 5058 752 5110 808
rect 4820 728 5110 752
rect 4820 706 5002 728
rect 4820 654 4834 706
rect 4886 672 5002 706
rect 5058 672 5110 728
rect 4886 654 5110 672
rect 4820 648 5110 654
rect 4820 592 5002 648
rect 5058 592 5110 648
rect 4820 568 5110 592
rect 4820 512 5002 568
rect 5058 512 5110 568
rect 4820 506 5110 512
rect 4820 454 4834 506
rect 4886 488 5110 506
rect 4886 454 5002 488
rect 4820 432 5002 454
rect 5058 432 5110 488
rect 4820 408 5110 432
rect 4820 352 5002 408
rect 5058 352 5110 408
rect 4820 328 5110 352
rect 4820 316 5002 328
rect 4820 264 4834 316
rect 4886 272 5002 316
rect 5058 272 5110 328
rect 4886 264 5110 272
rect 4820 248 5110 264
rect 4820 192 5002 248
rect 5058 192 5110 248
rect 4820 168 5110 192
rect 4820 112 5002 168
rect 5058 112 5110 168
rect 4820 60 5110 112
rect 4520 -166 4714 -114
rect 4766 -166 4780 -114
rect 4520 -304 4780 -166
rect 4520 -356 4714 -304
rect 4766 -356 4780 -304
rect 4520 -724 4780 -356
rect 4820 -52 5110 10
rect 4820 -108 5002 -52
rect 5058 -108 5110 -52
rect 4820 -132 5110 -108
rect 4820 -188 5002 -132
rect 5058 -188 5110 -132
rect 4820 -204 5110 -188
rect 4820 -256 4834 -204
rect 4886 -212 5110 -204
rect 4886 -256 5002 -212
rect 4820 -268 5002 -256
rect 5058 -268 5110 -212
rect 4820 -292 5110 -268
rect 4820 -348 5002 -292
rect 5058 -348 5110 -292
rect 4820 -372 5110 -348
rect 4820 -394 5002 -372
rect 4820 -446 4834 -394
rect 4886 -428 5002 -394
rect 5058 -428 5110 -372
rect 4886 -446 5110 -428
rect 4820 -452 5110 -446
rect 4820 -508 5002 -452
rect 5058 -508 5110 -452
rect 4820 -550 5110 -508
rect 4820 -560 5080 -550
rect 4520 -776 4714 -724
rect 4766 -776 4780 -724
rect 4520 -914 4780 -776
rect 4520 -966 4714 -914
rect 4766 -966 4780 -914
rect 4520 -1150 4780 -966
rect 4820 -652 5110 -610
rect 4820 -708 5002 -652
rect 5058 -708 5110 -652
rect 4820 -732 5110 -708
rect 4820 -788 5002 -732
rect 5058 -788 5110 -732
rect 4820 -812 5110 -788
rect 4820 -824 5002 -812
rect 4820 -876 4834 -824
rect 4886 -868 5002 -824
rect 5058 -868 5110 -812
rect 4886 -876 5110 -868
rect 4820 -892 5110 -876
rect 4820 -948 5002 -892
rect 5058 -948 5110 -892
rect 4820 -972 5110 -948
rect 4820 -1028 5002 -972
rect 5058 -1028 5110 -972
rect 4820 -1060 5110 -1028
rect 4820 -1070 5080 -1060
rect 3730 -1217 3990 -1150
rect 3730 -1273 3792 -1217
rect 3848 -1254 3990 -1217
rect 3848 -1273 3924 -1254
rect 3730 -1297 3924 -1273
rect 3730 -1353 3792 -1297
rect 3848 -1306 3924 -1297
rect 3976 -1306 3990 -1254
rect 3848 -1353 3990 -1306
rect 3730 -1377 3990 -1353
rect 3730 -1433 3792 -1377
rect 3848 -1433 3990 -1377
rect 3730 -1510 3990 -1433
rect 4030 -1254 4780 -1150
rect 4030 -1294 4714 -1254
rect 4030 -1346 4347 -1294
rect 4399 -1346 4411 -1294
rect 4463 -1306 4714 -1294
rect 4766 -1306 4780 -1254
rect 4463 -1346 4780 -1306
rect 4030 -1354 4780 -1346
rect 4030 -1406 4044 -1354
rect 4096 -1406 4780 -1354
rect 4030 -1510 4780 -1406
rect 4820 -1182 5080 -1150
rect 4820 -1238 4972 -1182
rect 5028 -1238 5080 -1182
rect 4820 -1262 5080 -1238
rect 4820 -1318 4972 -1262
rect 5028 -1318 5080 -1262
rect 4820 -1342 5080 -1318
rect 4820 -1354 4972 -1342
rect 4820 -1406 4834 -1354
rect 4886 -1398 4972 -1354
rect 5028 -1398 5080 -1342
rect 4886 -1406 5080 -1398
rect 4820 -1422 5080 -1406
rect 4820 -1478 4972 -1422
rect 5028 -1478 5080 -1422
rect 4820 -1510 5080 -1478
<< via2 >>
rect 5002 832 5058 888
rect 5002 752 5058 808
rect 5002 672 5058 728
rect 5002 592 5058 648
rect 5002 512 5058 568
rect 5002 432 5058 488
rect 5002 352 5058 408
rect 5002 272 5058 328
rect 5002 192 5058 248
rect 5002 112 5058 168
rect 5002 -108 5058 -52
rect 5002 -188 5058 -132
rect 5002 -268 5058 -212
rect 5002 -348 5058 -292
rect 5002 -428 5058 -372
rect 5002 -508 5058 -452
rect 5002 -708 5058 -652
rect 5002 -788 5058 -732
rect 5002 -868 5058 -812
rect 5002 -948 5058 -892
rect 5002 -1028 5058 -972
rect 3792 -1273 3848 -1217
rect 3792 -1353 3848 -1297
rect 3792 -1433 3848 -1377
rect 4972 -1238 5028 -1182
rect 4972 -1318 5028 -1262
rect 4972 -1398 5028 -1342
rect 4972 -1478 5028 -1422
<< metal3 >>
rect 4950 892 5110 920
rect 4950 828 4998 892
rect 5062 828 5110 892
rect 4950 812 5110 828
rect 4950 748 4998 812
rect 5062 748 5110 812
rect 4950 732 5110 748
rect 4950 668 4998 732
rect 5062 668 5110 732
rect 4950 652 5110 668
rect 4950 588 4998 652
rect 5062 588 5110 652
rect 4950 572 5110 588
rect 4950 508 4998 572
rect 5062 508 5110 572
rect 4950 492 5110 508
rect 4950 428 4998 492
rect 5062 428 5110 492
rect 4950 412 5110 428
rect 4950 348 4998 412
rect 5062 348 5110 412
rect 4950 332 5110 348
rect 4950 268 4998 332
rect 5062 268 5110 332
rect 4950 252 5110 268
rect 4950 188 4998 252
rect 5062 188 5110 252
rect 4950 172 5110 188
rect 4950 108 4998 172
rect 5062 108 5110 172
rect 4950 60 5110 108
rect 4950 -48 5110 0
rect 4950 -112 4998 -48
rect 5062 -112 5110 -48
rect 4950 -128 5110 -112
rect 4950 -192 4998 -128
rect 5062 -192 5110 -128
rect 4950 -208 5110 -192
rect 4950 -272 4998 -208
rect 5062 -272 5110 -208
rect 4950 -288 5110 -272
rect 4950 -352 4998 -288
rect 5062 -352 5110 -288
rect 4950 -368 5110 -352
rect 4950 -432 4998 -368
rect 5062 -432 5110 -368
rect 4950 -448 5110 -432
rect 4950 -512 4998 -448
rect 5062 -512 5110 -448
rect 4950 -550 5110 -512
rect 4950 -652 5110 -630
rect 4950 -688 5002 -652
rect 5058 -688 5110 -652
rect 4950 -752 4998 -688
rect 5062 -752 5110 -688
rect 4950 -768 5002 -752
rect 5058 -768 5110 -752
rect 4950 -832 4998 -768
rect 5062 -832 5110 -768
rect 4950 -848 5002 -832
rect 5058 -848 5110 -832
rect 4950 -912 4998 -848
rect 5062 -912 5110 -848
rect 4950 -928 5002 -912
rect 5058 -928 5110 -912
rect 4950 -992 4998 -928
rect 5062 -992 5110 -928
rect 4950 -1028 5002 -992
rect 5058 -1028 5110 -992
rect 4950 -1060 5110 -1028
rect 3730 -1213 3900 -1150
rect 3730 -1277 3788 -1213
rect 3852 -1277 3900 -1213
rect 3730 -1293 3900 -1277
rect 3730 -1357 3788 -1293
rect 3852 -1357 3900 -1293
rect 3730 -1373 3900 -1357
rect 3730 -1437 3788 -1373
rect 3852 -1437 3900 -1373
rect 3730 -1510 3900 -1437
rect 4920 -1182 5080 -1150
rect 4920 -1218 4972 -1182
rect 5028 -1218 5080 -1182
rect 4920 -1282 4968 -1218
rect 5032 -1282 5080 -1218
rect 4920 -1298 4972 -1282
rect 5028 -1298 5080 -1282
rect 4920 -1362 4968 -1298
rect 5032 -1362 5080 -1298
rect 4920 -1378 4972 -1362
rect 5028 -1378 5080 -1362
rect 4920 -1442 4968 -1378
rect 5032 -1442 5080 -1378
rect 4920 -1478 4972 -1442
rect 5028 -1478 5080 -1442
rect 4920 -1510 5080 -1478
<< via3 >>
rect 4998 888 5062 892
rect 4998 832 5002 888
rect 5002 832 5058 888
rect 5058 832 5062 888
rect 4998 828 5062 832
rect 4998 808 5062 812
rect 4998 752 5002 808
rect 5002 752 5058 808
rect 5058 752 5062 808
rect 4998 748 5062 752
rect 4998 728 5062 732
rect 4998 672 5002 728
rect 5002 672 5058 728
rect 5058 672 5062 728
rect 4998 668 5062 672
rect 4998 648 5062 652
rect 4998 592 5002 648
rect 5002 592 5058 648
rect 5058 592 5062 648
rect 4998 588 5062 592
rect 4998 568 5062 572
rect 4998 512 5002 568
rect 5002 512 5058 568
rect 5058 512 5062 568
rect 4998 508 5062 512
rect 4998 488 5062 492
rect 4998 432 5002 488
rect 5002 432 5058 488
rect 5058 432 5062 488
rect 4998 428 5062 432
rect 4998 408 5062 412
rect 4998 352 5002 408
rect 5002 352 5058 408
rect 5058 352 5062 408
rect 4998 348 5062 352
rect 4998 328 5062 332
rect 4998 272 5002 328
rect 5002 272 5058 328
rect 5058 272 5062 328
rect 4998 268 5062 272
rect 4998 248 5062 252
rect 4998 192 5002 248
rect 5002 192 5058 248
rect 5058 192 5062 248
rect 4998 188 5062 192
rect 4998 168 5062 172
rect 4998 112 5002 168
rect 5002 112 5058 168
rect 5058 112 5062 168
rect 4998 108 5062 112
rect 4998 -52 5062 -48
rect 4998 -108 5002 -52
rect 5002 -108 5058 -52
rect 5058 -108 5062 -52
rect 4998 -112 5062 -108
rect 4998 -132 5062 -128
rect 4998 -188 5002 -132
rect 5002 -188 5058 -132
rect 5058 -188 5062 -132
rect 4998 -192 5062 -188
rect 4998 -212 5062 -208
rect 4998 -268 5002 -212
rect 5002 -268 5058 -212
rect 5058 -268 5062 -212
rect 4998 -272 5062 -268
rect 4998 -292 5062 -288
rect 4998 -348 5002 -292
rect 5002 -348 5058 -292
rect 5058 -348 5062 -292
rect 4998 -352 5062 -348
rect 4998 -372 5062 -368
rect 4998 -428 5002 -372
rect 5002 -428 5058 -372
rect 5058 -428 5062 -372
rect 4998 -432 5062 -428
rect 4998 -452 5062 -448
rect 4998 -508 5002 -452
rect 5002 -508 5058 -452
rect 5058 -508 5062 -452
rect 4998 -512 5062 -508
rect 4998 -708 5002 -688
rect 5002 -708 5058 -688
rect 5058 -708 5062 -688
rect 4998 -732 5062 -708
rect 4998 -752 5002 -732
rect 5002 -752 5058 -732
rect 5058 -752 5062 -732
rect 4998 -788 5002 -768
rect 5002 -788 5058 -768
rect 5058 -788 5062 -768
rect 4998 -812 5062 -788
rect 4998 -832 5002 -812
rect 5002 -832 5058 -812
rect 5058 -832 5062 -812
rect 4998 -868 5002 -848
rect 5002 -868 5058 -848
rect 5058 -868 5062 -848
rect 4998 -892 5062 -868
rect 4998 -912 5002 -892
rect 5002 -912 5058 -892
rect 5058 -912 5062 -892
rect 4998 -948 5002 -928
rect 5002 -948 5058 -928
rect 5058 -948 5062 -928
rect 4998 -972 5062 -948
rect 4998 -992 5002 -972
rect 5002 -992 5058 -972
rect 5058 -992 5062 -972
rect 3788 -1217 3852 -1213
rect 3788 -1273 3792 -1217
rect 3792 -1273 3848 -1217
rect 3848 -1273 3852 -1217
rect 3788 -1277 3852 -1273
rect 3788 -1297 3852 -1293
rect 3788 -1353 3792 -1297
rect 3792 -1353 3848 -1297
rect 3848 -1353 3852 -1297
rect 3788 -1357 3852 -1353
rect 3788 -1377 3852 -1373
rect 3788 -1433 3792 -1377
rect 3792 -1433 3848 -1377
rect 3848 -1433 3852 -1377
rect 3788 -1437 3852 -1433
rect 4968 -1238 4972 -1218
rect 4972 -1238 5028 -1218
rect 5028 -1238 5032 -1218
rect 4968 -1262 5032 -1238
rect 4968 -1282 4972 -1262
rect 4972 -1282 5028 -1262
rect 5028 -1282 5032 -1262
rect 4968 -1318 4972 -1298
rect 4972 -1318 5028 -1298
rect 5028 -1318 5032 -1298
rect 4968 -1342 5032 -1318
rect 4968 -1362 4972 -1342
rect 4972 -1362 5028 -1342
rect 5028 -1362 5032 -1342
rect 4968 -1398 4972 -1378
rect 4972 -1398 5028 -1378
rect 5028 -1398 5032 -1378
rect 4968 -1422 5032 -1398
rect 4968 -1442 4972 -1422
rect 4972 -1442 5028 -1422
rect 5028 -1442 5032 -1422
<< metal4 >>
rect 4370 2260 4890 2540
rect 3730 -1213 4090 -500
rect 4510 -630 4670 1930
rect 4730 0 4890 2260
rect 4950 892 5110 4368
rect 4950 828 4998 892
rect 5062 828 5110 892
rect 4950 812 5110 828
rect 4950 748 4998 812
rect 5062 748 5110 812
rect 4950 732 5110 748
rect 4950 668 4998 732
rect 5062 668 5110 732
rect 4950 652 5110 668
rect 4950 588 4998 652
rect 5062 588 5110 652
rect 4950 572 5110 588
rect 4950 508 4998 572
rect 5062 508 5110 572
rect 4950 492 5110 508
rect 4950 428 4998 492
rect 5062 428 5110 492
rect 4950 412 5110 428
rect 4950 348 4998 412
rect 5062 348 5110 412
rect 4950 332 5110 348
rect 4950 268 4998 332
rect 5062 268 5110 332
rect 4950 252 5110 268
rect 4950 188 4998 252
rect 5062 188 5110 252
rect 4950 172 5110 188
rect 4950 108 4998 172
rect 5062 108 5110 172
rect 4950 60 5110 108
rect 4730 -48 5110 0
rect 4730 -112 4998 -48
rect 5062 -112 5110 -48
rect 4730 -128 5110 -112
rect 4730 -192 4998 -128
rect 5062 -192 5110 -128
rect 4730 -208 5110 -192
rect 4730 -272 4998 -208
rect 5062 -272 5110 -208
rect 4730 -288 5110 -272
rect 4730 -352 4998 -288
rect 5062 -352 5110 -288
rect 4730 -368 5110 -352
rect 4730 -432 4998 -368
rect 5062 -432 5110 -368
rect 4730 -448 5110 -432
rect 4730 -512 4998 -448
rect 5062 -512 5110 -448
rect 4730 -560 5110 -512
rect 4510 -688 5110 -630
rect 4510 -752 4998 -688
rect 5062 -752 5110 -688
rect 4510 -768 5110 -752
rect 4510 -832 4998 -768
rect 5062 -832 5110 -768
rect 4510 -848 5110 -832
rect 4510 -912 4998 -848
rect 5062 -912 5110 -848
rect 4510 -928 5110 -912
rect 4510 -992 4998 -928
rect 5062 -992 5110 -928
rect 4510 -1060 5110 -992
rect 4510 -1070 5080 -1060
rect 3730 -1277 3788 -1213
rect 3852 -1277 4090 -1213
rect 3730 -1293 4090 -1277
rect 3730 -1357 3788 -1293
rect 3852 -1357 4090 -1293
rect 3730 -1373 4090 -1357
rect 3730 -1437 3788 -1373
rect 3852 -1437 4090 -1373
rect 3730 -1510 4090 -1437
rect 4760 -1212 5080 -1150
rect 4760 -1448 4812 -1212
rect 5048 -1448 5080 -1212
rect 4760 -1510 5080 -1448
<< via4 >>
rect 4812 -1218 5048 -1212
rect 4812 -1282 4968 -1218
rect 4968 -1282 5032 -1218
rect 5032 -1282 5048 -1218
rect 4812 -1298 5048 -1282
rect 4812 -1362 4968 -1298
rect 4968 -1362 5032 -1298
rect 5032 -1362 5048 -1298
rect 4812 -1378 5048 -1362
rect 4812 -1442 4968 -1378
rect 4968 -1442 5032 -1378
rect 5032 -1442 5048 -1378
rect 4812 -1448 5048 -1442
<< metal5 >>
rect 3380 3710 4990 4830
rect 3380 3700 4930 3710
rect 3380 1430 3970 3700
rect 3380 -420 3780 1430
rect 4280 400 5080 1000
rect 4760 -1212 5080 400
rect 4760 -1448 4812 -1212
rect 5048 -1448 5080 -1212
rect 4760 -1510 5080 -1448
use sky130_fd_pr__cap_mim_m3_2_WCTBV5  XC1
timestamp 1663011646
transform 1 0 3851 0 1 701
box -551 -301 573 301
use sky130_fd_pr__cap_mim_m3_2_WCTZRP  XC2
timestamp 1663011646
transform 1 0 3951 0 1 1631
box -651 -301 673 301
use sky130_fd_pr__cap_mim_m3_2_3ZFDVT  XC3
timestamp 1663011646
transform 1 0 3951 0 1 2761
box -651 -501 673 501
use sky130_fd_pr__cap_mim_m3_2_VCH7EQ  XC4
timestamp 1663011646
transform 0 1 4611 1 0 4541
box -951 -501 973 501
use sky130_fd_pr__cap_mim_m3_2_FJFAMD  XC6
timestamp 1663011646
transform 1 0 3851 0 1 -229
box -551 -301 573 301
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM1
timestamp 1663011646
transform 0 1 4010 -1 0 -1329
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM2
timestamp 1663011646
transform 0 1 4800 -1 0 -1329
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_lvt_DJ7QE5  XM3
timestamp 1663011646
transform 0 -1 4800 1 0 -847
box -253 -300 253 300
use sky130_fd_pr__nfet_01v8_lvt_BX7S53  XM4
timestamp 1663011646
transform 0 1 4800 -1 0 -279
box -301 -300 301 300
use sky130_fd_pr__nfet_01v8_lvt_B6HS5D  XM5
timestamp 1663011646
transform 0 1 4800 -1 0 485
box -445 -300 445 300
<< labels >>
rlabel metal2 s 4100 -1510 4710 -1150 4 GND
port 1 nsew
rlabel metal5 s 3380 3700 4930 4830 4 IN
port 2 nsew
rlabel metal1 s 3300 -1540 5110 -1480 4 ctrll1
port 3 nsew
rlabel metal1 s 3300 -1180 5110 -1120 4 ctrll2
port 4 nsew
rlabel metal1 s 3300 -640 5110 -580 4 ctrll3
port 5 nsew
rlabel metal1 s 3300 -50 5110 10 4 ctrll4
port 6 nsew
rlabel metal1 s 3300 860 5110 920 4 ctrll5
port 7 nsew
<< end >>
