magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 6405 3125 6675 3160
rect 7100 3125 7370 3160
rect 7840 3125 8110 3160
rect 6410 1935 6680 1970
rect 7135 1935 7405 1970
rect 7840 1935 8110 1970
rect 6410 1750 6680 1785
rect 7145 1750 7415 1785
rect 7830 1750 8100 1785
rect 6405 1435 6675 1470
rect 7145 1435 7415 1470
rect 7850 1435 8120 1470
<< metal1 >>
rect 5155 8478 6315 8510
rect 5155 8106 5197 8478
rect 6273 8106 6315 8478
rect 5155 8075 6315 8106
rect 8200 8478 9360 8510
rect 8200 8106 8242 8478
rect 9318 8106 9360 8478
rect 8200 8075 9360 8106
rect 5000 3125 9520 3185
rect 6720 2085 6780 3125
rect 6810 3050 6895 3060
rect 6810 3048 7010 3050
rect 6810 2996 6826 3048
rect 6878 3000 7010 3048
rect 6878 2996 6895 3000
rect 6810 2990 6895 2996
rect 6930 2963 7010 2970
rect 6930 2956 6944 2963
rect 6810 2911 6944 2956
rect 6996 2911 7010 2963
rect 6810 2905 7010 2911
rect 6930 2900 7010 2905
rect 6810 2863 6895 2875
rect 6810 2811 6826 2863
rect 6878 2860 6895 2863
rect 6878 2811 7010 2860
rect 6810 2810 7010 2811
rect 6810 2805 6895 2810
rect 6930 2768 7010 2780
rect 6930 2762 6944 2768
rect 6810 2716 6944 2762
rect 6996 2716 7010 2768
rect 6810 2710 7010 2716
rect 6930 2705 7010 2710
rect 6810 2670 6895 2680
rect 6810 2668 7010 2670
rect 6810 2616 6826 2668
rect 6878 2620 7010 2668
rect 6878 2616 6895 2620
rect 6810 2605 6895 2616
rect 6930 2578 7010 2590
rect 6930 2571 6944 2578
rect 6810 2526 6944 2571
rect 6996 2526 7010 2578
rect 6810 2520 7010 2526
rect 6930 2515 7010 2520
rect 6810 2478 6895 2490
rect 6810 2426 6826 2478
rect 6878 2475 6895 2478
rect 6878 2426 7010 2475
rect 6810 2425 7010 2426
rect 6810 2415 6895 2425
rect 6930 2383 7010 2395
rect 6930 2378 6944 2383
rect 6810 2331 6944 2378
rect 6996 2331 7010 2383
rect 6810 2325 7010 2331
rect 6930 2320 7010 2325
rect 6810 2285 6895 2295
rect 6810 2283 7010 2285
rect 6810 2231 6826 2283
rect 6878 2235 7010 2283
rect 6878 2231 6895 2235
rect 6810 2220 6895 2231
rect 6930 2193 7010 2205
rect 6930 2186 6944 2193
rect 6810 2141 6944 2186
rect 6996 2141 7010 2193
rect 7040 2175 7100 3125
rect 7420 2175 7480 3125
rect 7625 3050 7710 3060
rect 7510 3048 7710 3050
rect 7510 3000 7641 3048
rect 7625 2996 7641 3000
rect 7693 2996 7710 3048
rect 7625 2990 7710 2996
rect 7510 2963 7590 2970
rect 7510 2911 7524 2963
rect 7576 2956 7590 2963
rect 7576 2911 7710 2956
rect 7510 2905 7710 2911
rect 7510 2900 7590 2905
rect 7625 2863 7710 2875
rect 7625 2860 7641 2863
rect 7510 2811 7641 2860
rect 7693 2811 7710 2863
rect 7510 2810 7710 2811
rect 7625 2805 7710 2810
rect 7510 2768 7590 2780
rect 7510 2716 7524 2768
rect 7576 2761 7590 2768
rect 7576 2716 7710 2761
rect 7510 2710 7710 2716
rect 7510 2705 7590 2710
rect 7625 2670 7710 2680
rect 7510 2668 7710 2670
rect 7510 2620 7641 2668
rect 7625 2616 7641 2620
rect 7693 2616 7710 2668
rect 7625 2605 7710 2616
rect 7510 2578 7590 2590
rect 7510 2526 7524 2578
rect 7576 2571 7590 2578
rect 7576 2526 7710 2571
rect 7510 2520 7710 2526
rect 7510 2515 7590 2520
rect 7625 2478 7710 2490
rect 7625 2475 7641 2478
rect 7510 2426 7641 2475
rect 7693 2426 7710 2478
rect 7510 2425 7710 2426
rect 7625 2415 7710 2425
rect 7510 2383 7590 2390
rect 7510 2331 7524 2383
rect 7576 2376 7590 2383
rect 7576 2331 7710 2376
rect 7510 2325 7710 2331
rect 7510 2320 7590 2325
rect 7625 2285 7710 2295
rect 7510 2283 7710 2285
rect 7510 2235 7641 2283
rect 7625 2231 7641 2235
rect 7693 2231 7710 2283
rect 7625 2220 7710 2231
rect 7510 2193 7590 2205
rect 6810 2135 7010 2141
rect 6930 2130 7010 2135
rect 7510 2141 7524 2193
rect 7576 2185 7590 2193
rect 7576 2141 7710 2185
rect 7510 2135 7710 2141
rect 7510 2130 7590 2135
rect 6810 2093 6895 2105
rect 6810 2041 6826 2093
rect 6878 2090 6895 2093
rect 7625 2093 7710 2105
rect 7625 2090 7641 2093
rect 6878 2041 7015 2090
rect 6810 2040 7015 2041
rect 7505 2041 7641 2090
rect 7693 2041 7710 2093
rect 7740 2085 7800 3125
rect 7505 2040 7710 2041
rect 6810 2035 6895 2040
rect 7625 2035 7710 2040
rect 5165 1968 6315 2000
rect 5165 1596 5202 1968
rect 6278 1596 6315 1968
rect 8205 1968 9350 1995
rect 6810 1703 7010 1725
rect 6810 1651 6820 1703
rect 6872 1651 6884 1703
rect 6936 1651 6948 1703
rect 7000 1651 7010 1703
rect 5165 1565 6315 1596
rect 6730 1450 6780 1645
rect 6810 1630 7010 1651
rect 7510 1703 7710 1725
rect 7510 1651 7520 1703
rect 7572 1651 7584 1703
rect 7636 1651 7648 1703
rect 7700 1651 7710 1703
rect 6810 1573 7010 1590
rect 6810 1521 6820 1573
rect 6872 1521 6884 1573
rect 6936 1521 6948 1573
rect 7000 1521 7010 1573
rect 6810 1505 7010 1521
rect 7040 1450 7090 1645
rect 6730 1400 7090 1450
rect 7430 1450 7480 1645
rect 7510 1630 7710 1651
rect 7510 1573 7710 1590
rect 7510 1521 7520 1573
rect 7572 1521 7584 1573
rect 7636 1521 7648 1573
rect 7700 1521 7710 1573
rect 7510 1505 7710 1521
rect 7740 1450 7790 1645
rect 8205 1596 8242 1968
rect 9318 1596 9350 1968
rect 8205 1565 9350 1596
rect 7430 1400 7790 1450
<< via1 >>
rect 5197 8106 6273 8478
rect 8242 8106 9318 8478
rect 6826 2996 6878 3048
rect 6944 2911 6996 2963
rect 6826 2811 6878 2863
rect 6944 2716 6996 2768
rect 6826 2616 6878 2668
rect 6944 2526 6996 2578
rect 6826 2426 6878 2478
rect 6944 2331 6996 2383
rect 6826 2231 6878 2283
rect 6944 2141 6996 2193
rect 7641 2996 7693 3048
rect 7524 2911 7576 2963
rect 7641 2811 7693 2863
rect 7524 2716 7576 2768
rect 7641 2616 7693 2668
rect 7524 2526 7576 2578
rect 7641 2426 7693 2478
rect 7524 2331 7576 2383
rect 7641 2231 7693 2283
rect 7524 2141 7576 2193
rect 6826 2041 6878 2093
rect 7641 2041 7693 2093
rect 5202 1596 6278 1968
rect 6820 1651 6872 1703
rect 6884 1651 6936 1703
rect 6948 1651 7000 1703
rect 7520 1651 7572 1703
rect 7584 1651 7636 1703
rect 7648 1651 7700 1703
rect 6820 1521 6872 1573
rect 6884 1521 6936 1573
rect 6948 1521 7000 1573
rect 7520 1521 7572 1573
rect 7584 1521 7636 1573
rect 7648 1521 7700 1573
rect 8242 1596 9318 1968
<< metal2 >>
rect 5000 8478 9520 8510
rect 5000 8106 5197 8478
rect 6273 8106 8242 8478
rect 9318 8106 9520 8478
rect 5000 8070 9520 8106
rect 5000 3225 9520 3625
rect 6495 3048 6895 3225
rect 6495 2996 6826 3048
rect 6878 2996 6895 3048
rect 6495 2863 6895 2996
rect 7040 2975 7480 3065
rect 7625 3048 8025 3225
rect 7625 2996 7641 3048
rect 7693 2996 8025 3048
rect 6930 2963 7590 2975
rect 6930 2911 6944 2963
rect 6996 2911 7524 2963
rect 7576 2911 7590 2963
rect 6930 2900 7590 2911
rect 6495 2811 6826 2863
rect 6878 2811 6895 2863
rect 6495 2668 6895 2811
rect 7040 2780 7480 2900
rect 7625 2863 8025 2996
rect 7625 2811 7641 2863
rect 7693 2811 8025 2863
rect 6930 2768 7590 2780
rect 6930 2716 6944 2768
rect 6996 2716 7524 2768
rect 7576 2716 7590 2768
rect 6930 2705 7590 2716
rect 6495 2616 6826 2668
rect 6878 2616 6895 2668
rect 6495 2478 6895 2616
rect 7040 2590 7480 2705
rect 7625 2668 8025 2811
rect 7625 2616 7641 2668
rect 7693 2616 8025 2668
rect 6930 2578 7590 2590
rect 6930 2526 6944 2578
rect 6996 2526 7524 2578
rect 7576 2526 7590 2578
rect 6930 2515 7590 2526
rect 6495 2426 6826 2478
rect 6878 2426 6895 2478
rect 6495 2283 6895 2426
rect 7040 2395 7480 2515
rect 7625 2478 8025 2616
rect 7625 2426 7641 2478
rect 7693 2426 8025 2478
rect 6930 2383 7590 2395
rect 6930 2331 6944 2383
rect 6996 2331 7524 2383
rect 7576 2331 7590 2383
rect 6930 2320 7590 2331
rect 6495 2231 6826 2283
rect 6878 2231 6895 2283
rect 6495 2093 6895 2231
rect 7040 2205 7480 2320
rect 7625 2283 8025 2426
rect 7625 2231 7641 2283
rect 7693 2231 8025 2283
rect 6930 2193 7590 2205
rect 6930 2141 6944 2193
rect 6996 2141 7524 2193
rect 7576 2141 7590 2193
rect 6930 2130 7590 2141
rect 6495 2041 6826 2093
rect 6878 2041 6895 2093
rect 6495 2035 6895 2041
rect 5165 1970 6315 2000
rect 5165 1594 5192 1970
rect 6288 1594 6315 1970
rect 7040 1870 7480 2130
rect 7625 2093 8025 2231
rect 7625 2041 7641 2093
rect 7693 2041 8025 2093
rect 7625 2035 8025 2041
rect 8205 1970 9350 2000
rect 6715 1720 7805 1870
rect 6715 1703 7105 1720
rect 6715 1685 6820 1703
rect 6810 1651 6820 1685
rect 6872 1651 6884 1703
rect 6936 1651 6948 1703
rect 7000 1685 7105 1703
rect 7415 1703 7805 1720
rect 7415 1685 7520 1703
rect 7000 1651 7010 1685
rect 6810 1630 7010 1651
rect 7510 1651 7520 1685
rect 7572 1651 7584 1703
rect 7636 1651 7648 1703
rect 7700 1685 7805 1703
rect 7700 1651 7710 1685
rect 7510 1630 7710 1651
rect 5165 1565 6315 1594
rect 8205 1594 8232 1970
rect 9328 1594 9350 1970
rect 6810 1575 7010 1590
rect 6810 1573 6842 1575
rect 6898 1573 6922 1575
rect 6978 1573 7010 1575
rect 6810 1521 6820 1573
rect 7000 1521 7010 1573
rect 6810 1519 6842 1521
rect 6898 1519 6922 1521
rect 6978 1519 7010 1521
rect 6810 1505 7010 1519
rect 7510 1575 7710 1590
rect 7510 1573 7542 1575
rect 7598 1573 7622 1575
rect 7678 1573 7710 1575
rect 7510 1521 7520 1573
rect 7700 1521 7710 1573
rect 8205 1570 9350 1594
rect 7510 1519 7542 1521
rect 7598 1519 7622 1521
rect 7678 1519 7710 1521
rect 7510 1505 7710 1519
<< via2 >>
rect 5192 1968 6288 1970
rect 5192 1596 5202 1968
rect 5202 1596 6278 1968
rect 6278 1596 6288 1968
rect 5192 1594 6288 1596
rect 8232 1968 9328 1970
rect 8232 1596 8242 1968
rect 8242 1596 9318 1968
rect 9318 1596 9328 1968
rect 8232 1594 9328 1596
rect 6842 1573 6898 1575
rect 6922 1573 6978 1575
rect 6842 1521 6872 1573
rect 6872 1521 6884 1573
rect 6884 1521 6898 1573
rect 6922 1521 6936 1573
rect 6936 1521 6948 1573
rect 6948 1521 6978 1573
rect 6842 1519 6898 1521
rect 6922 1519 6978 1521
rect 7542 1573 7598 1575
rect 7622 1573 7678 1575
rect 7542 1521 7572 1573
rect 7572 1521 7584 1573
rect 7584 1521 7598 1573
rect 7622 1521 7636 1573
rect 7636 1521 7648 1573
rect 7648 1521 7678 1573
rect 7542 1519 7598 1521
rect 7622 1519 7678 1521
<< metal3 >>
rect 5165 1970 6315 2000
rect 5165 1594 5192 1970
rect 6288 1594 6315 1970
rect 5165 1590 6315 1594
rect 8205 1970 9350 1995
rect 8205 1594 8232 1970
rect 9328 1594 9350 1970
rect 8205 1590 9350 1594
rect 5165 1575 7010 1590
rect 5165 1519 6842 1575
rect 6898 1519 6922 1575
rect 6978 1519 7010 1575
rect 5165 1410 7010 1519
rect 7510 1575 9350 1590
rect 7510 1519 7542 1575
rect 7598 1519 7622 1575
rect 7678 1519 9350 1575
rect 7510 1410 9350 1519
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM1
timestamp 1663011646
transform 0 -1 6910 -1 0 2547
box -637 -300 637 300
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM2
timestamp 1663011646
transform 0 1 6910 -1 0 1611
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_lvt_648S5X  XM3
timestamp 1663011646
transform 0 1 7610 -1 0 1611
box -201 -300 201 300
use sky130_fd_pr__nfet_01v8_lvt_9DHFGX  XM4
timestamp 1663011646
transform 0 1 7610 -1 0 2547
box -637 -300 637 300
use sky130_fd_pr__res_high_po_5p73_YZEQ6M  XR1
timestamp 1663011646
transform 1 0 5739 0 1 5038
box -729 -3628 729 3628
use sky130_fd_pr__res_high_po_5p73_YZEQ6M  XR2
timestamp 1663011646
transform 1 0 8779 0 1 5038
box -729 -3628 729 3628
<< labels >>
rlabel metal1 s 7430 1400 7790 1450 4 INA
port 1 nsew
rlabel metal1 s 6730 1400 7090 1450 4 INB
port 2 nsew
rlabel metal1 s 5000 3125 9520 3185 4 BIAS
port 3 nsew
rlabel metal2 s 5000 3225 9520 3625 4 GND
port 4 nsew
rlabel metal2 s 6295 8075 8220 8510 4 VDD
port 5 nsew
rlabel metal3 s 5165 1410 6820 1585 4 OUTB
port 6 nsew
rlabel metal3 s 7700 1410 9350 1585 4 OUTA
port 7 nsew
rlabel locali s 7145 1435 7415 1470 4 SUB
port 8 nsew
<< end >>
