magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -140 -160 2080 1600
<< nsubdiff >>
rect -60 1557 2000 1560
rect -60 1523 885 1557
rect 919 1523 953 1557
rect 987 1523 1021 1557
rect 1055 1523 2000 1557
rect -60 1520 2000 1523
rect -60 859 -20 1520
rect -60 825 -57 859
rect -23 825 -20 859
rect -60 791 -20 825
rect -60 757 -57 791
rect -23 757 -20 791
rect -60 723 -20 757
rect -60 689 -57 723
rect -23 689 -20 723
rect -60 655 -20 689
rect -60 621 -57 655
rect -23 621 -20 655
rect -60 -40 -20 621
rect 1960 859 2000 1520
rect 1960 825 1963 859
rect 1997 825 2000 859
rect 1960 791 2000 825
rect 1960 757 1963 791
rect 1997 757 2000 791
rect 1960 723 2000 757
rect 1960 689 1963 723
rect 1997 689 2000 723
rect 1960 655 2000 689
rect 1960 621 1963 655
rect 1997 621 2000 655
rect 1960 -40 2000 621
rect -60 -43 2000 -40
rect -60 -77 885 -43
rect 919 -77 953 -43
rect 987 -77 1021 -43
rect 1055 -77 2000 -43
rect -60 -80 2000 -77
<< nsubdiffcont >>
rect 885 1523 919 1557
rect 953 1523 987 1557
rect 1021 1523 1055 1557
rect -57 825 -23 859
rect -57 757 -23 791
rect -57 689 -23 723
rect -57 621 -23 655
rect 1963 825 1997 859
rect 1963 757 1997 791
rect 1963 689 1997 723
rect 1963 621 1997 655
rect 885 -77 919 -43
rect 953 -77 987 -43
rect 1021 -77 1055 -43
<< locali >>
rect -60 1557 2000 1560
rect -60 1523 885 1557
rect 919 1523 953 1557
rect 987 1523 1021 1557
rect 1055 1523 2000 1557
rect -60 1520 2000 1523
rect -60 859 -20 1520
rect -60 825 -57 859
rect -23 825 -20 859
rect -60 791 -20 825
rect -60 757 -57 791
rect -23 757 -20 791
rect -60 723 -20 757
rect -60 689 -57 723
rect -23 689 -20 723
rect -60 655 -20 689
rect -60 621 -57 655
rect -23 621 -20 655
rect -60 -40 -20 621
rect 1960 859 2000 1520
rect 1960 825 1963 859
rect 1997 825 2000 859
rect 1960 791 2000 825
rect 1960 757 1963 791
rect 1997 757 2000 791
rect 1960 723 2000 757
rect 1960 689 1963 723
rect 1997 689 2000 723
rect 1960 655 2000 689
rect 1960 621 1963 655
rect 1997 621 2000 655
rect 1960 -40 2000 621
rect -60 -43 2000 -40
rect -60 -77 885 -43
rect 919 -77 953 -43
rect 987 -77 1021 -43
rect 1055 -77 2000 -43
rect -60 -80 2000 -77
<< metal1 >>
rect 30 1396 110 1400
rect 30 1344 44 1396
rect 96 1344 110 1396
rect 30 1340 110 1344
rect 550 1396 630 1400
rect 550 1344 564 1396
rect 616 1344 630 1396
rect 550 1340 630 1344
rect 1070 1396 1150 1400
rect 1070 1344 1084 1396
rect 1136 1344 1150 1396
rect 1070 1340 1150 1344
rect 1570 1396 1650 1400
rect 1570 1344 1584 1396
rect 1636 1344 1650 1396
rect 1570 1340 1650 1344
rect 290 1256 370 1260
rect 290 1204 304 1256
rect 356 1204 370 1256
rect 290 1200 370 1204
rect 810 1256 890 1260
rect 810 1204 824 1256
rect 876 1204 890 1256
rect 810 1200 890 1204
rect 1330 1256 1410 1260
rect 1330 1204 1344 1256
rect 1396 1204 1410 1256
rect 1330 1200 1410 1204
rect 1830 1256 1910 1260
rect 1830 1204 1844 1256
rect 1896 1204 1910 1256
rect 1830 1200 1910 1204
rect 104 1108 1842 1154
rect 30 1036 110 1040
rect 30 984 44 1036
rect 96 984 110 1036
rect 30 980 110 984
rect 550 1036 630 1040
rect 550 984 564 1036
rect 616 984 630 1036
rect 550 980 630 984
rect 1070 1036 1150 1040
rect 1070 984 1084 1036
rect 1136 984 1150 1036
rect 1070 980 1150 984
rect 1570 1036 1650 1040
rect 1570 984 1584 1036
rect 1636 984 1650 1036
rect 1570 980 1650 984
rect 290 876 370 880
rect 290 824 304 876
rect 356 824 370 876
rect 290 820 370 824
rect 810 876 890 880
rect 810 824 824 876
rect 876 824 890 876
rect 810 820 890 824
rect 1310 876 1390 880
rect 1310 824 1324 876
rect 1376 824 1390 876
rect 1310 820 1390 824
rect 1830 876 1910 880
rect 1830 824 1844 876
rect 1896 824 1910 876
rect 1830 820 1910 824
rect 102 742 1840 788
rect 30 656 110 660
rect 30 604 44 656
rect 96 604 110 656
rect 30 600 110 604
rect 550 656 630 660
rect 550 604 564 656
rect 616 604 630 656
rect 550 600 630 604
rect 1050 656 1130 660
rect 1050 604 1064 656
rect 1116 604 1130 656
rect 1050 600 1130 604
rect 1570 656 1650 660
rect 1570 604 1584 656
rect 1636 604 1650 656
rect 1570 600 1650 604
rect 290 516 370 520
rect 290 464 304 516
rect 356 464 370 516
rect 290 460 370 464
rect 790 516 870 520
rect 790 464 804 516
rect 856 464 870 516
rect 790 460 870 464
rect 1310 516 1390 520
rect 1310 464 1324 516
rect 1376 464 1390 516
rect 1310 460 1390 464
rect 1830 516 1910 520
rect 1830 464 1844 516
rect 1896 464 1910 516
rect 1830 460 1910 464
rect 100 382 1838 428
rect 30 296 110 300
rect 30 244 44 296
rect 96 244 110 296
rect 30 240 110 244
rect 550 296 630 300
rect 550 244 564 296
rect 616 244 630 296
rect 550 240 630 244
rect 1050 296 1130 300
rect 1050 244 1064 296
rect 1116 244 1130 296
rect 1050 240 1130 244
rect 1570 296 1650 300
rect 1570 244 1584 296
rect 1636 244 1650 296
rect 1570 240 1650 244
rect 290 156 370 160
rect 290 104 304 156
rect 356 104 370 156
rect 290 100 370 104
rect 790 156 870 160
rect 790 104 804 156
rect 856 104 870 156
rect 790 100 870 104
rect 1310 156 1390 160
rect 1310 104 1324 156
rect 1376 104 1390 156
rect 1310 100 1390 104
rect 1830 156 1910 160
rect 1830 104 1844 156
rect 1896 104 1910 156
rect 1830 100 1910 104
rect 102 14 1840 60
<< via1 >>
rect 44 1344 96 1396
rect 564 1344 616 1396
rect 1084 1344 1136 1396
rect 1584 1344 1636 1396
rect 304 1204 356 1256
rect 824 1204 876 1256
rect 1344 1204 1396 1256
rect 1844 1204 1896 1256
rect 44 984 96 1036
rect 564 984 616 1036
rect 1084 984 1136 1036
rect 1584 984 1636 1036
rect 304 824 356 876
rect 824 824 876 876
rect 1324 824 1376 876
rect 1844 824 1896 876
rect 44 604 96 656
rect 564 604 616 656
rect 1064 604 1116 656
rect 1584 604 1636 656
rect 304 464 356 516
rect 804 464 856 516
rect 1324 464 1376 516
rect 1844 464 1896 516
rect 44 244 96 296
rect 564 244 616 296
rect 1064 244 1116 296
rect 1584 244 1636 296
rect 304 104 356 156
rect 804 104 856 156
rect 1324 104 1376 156
rect 1844 104 1896 156
<< metal2 >>
rect 40 1400 100 1410
rect 560 1400 620 1410
rect 1080 1400 1140 1410
rect 1580 1400 1640 1410
rect 40 1396 1640 1400
rect 40 1344 44 1396
rect 96 1344 564 1396
rect 616 1344 1084 1396
rect 1136 1344 1584 1396
rect 1636 1344 1640 1396
rect 40 1340 1640 1344
rect 40 1040 100 1340
rect 560 1330 620 1340
rect 1080 1330 1140 1340
rect 1580 1330 1640 1340
rect 300 1260 360 1270
rect 820 1260 880 1270
rect 1340 1260 1400 1270
rect 1840 1260 1900 1270
rect 300 1256 1900 1260
rect 300 1204 304 1256
rect 356 1204 824 1256
rect 876 1204 1344 1256
rect 1396 1204 1844 1256
rect 1896 1204 1900 1256
rect 300 1200 1900 1204
rect 300 1190 360 1200
rect 820 1190 880 1200
rect 1340 1190 1400 1200
rect 560 1040 620 1050
rect 1080 1040 1140 1050
rect 1580 1040 1640 1050
rect 40 1036 1640 1040
rect 40 984 44 1036
rect 96 984 564 1036
rect 616 984 1084 1036
rect 1136 984 1584 1036
rect 1636 984 1640 1036
rect 40 980 1640 984
rect 40 660 100 980
rect 560 970 620 980
rect 1080 970 1140 980
rect 1580 970 1640 980
rect 300 880 360 890
rect 820 880 880 890
rect 1320 880 1380 890
rect 1840 880 1900 1200
rect 300 876 1900 880
rect 300 824 304 876
rect 356 824 824 876
rect 876 824 1324 876
rect 1376 824 1844 876
rect 1896 824 1900 876
rect 300 820 1900 824
rect 300 810 360 820
rect 820 810 880 820
rect 1320 810 1380 820
rect 560 660 620 670
rect 1060 660 1120 670
rect 1580 660 1640 670
rect 40 656 1640 660
rect 40 604 44 656
rect 96 604 564 656
rect 616 604 1064 656
rect 1116 604 1584 656
rect 1636 604 1640 656
rect 40 600 1640 604
rect 40 300 100 600
rect 560 590 620 600
rect 1060 590 1120 600
rect 1580 590 1640 600
rect 300 520 360 530
rect 800 520 860 530
rect 1320 520 1380 530
rect 1840 520 1900 820
rect 300 516 1900 520
rect 300 464 304 516
rect 356 464 804 516
rect 856 464 1324 516
rect 1376 464 1844 516
rect 1896 464 1900 516
rect 300 460 1900 464
rect 300 450 360 460
rect 800 450 860 460
rect 1320 450 1380 460
rect 560 300 620 310
rect 1060 300 1120 310
rect 1580 300 1640 310
rect 40 296 1640 300
rect 40 244 44 296
rect 96 244 564 296
rect 616 244 1064 296
rect 1116 244 1584 296
rect 1636 244 1640 296
rect 40 240 1640 244
rect 40 230 100 240
rect 560 230 620 240
rect 1060 230 1120 240
rect 1580 230 1640 240
rect 300 160 360 170
rect 800 160 860 170
rect 1320 160 1380 170
rect 1840 160 1900 460
rect 300 156 1900 160
rect 300 104 304 156
rect 356 104 804 156
rect 856 104 1324 156
rect 1376 104 1844 156
rect 1896 104 1900 156
rect 300 100 1900 104
rect 300 90 360 100
rect 800 90 860 100
rect 1320 90 1380 100
rect 1840 90 1900 100
use sky130_fd_pr__pfet_01v8_lvt_9UM225  sky130_fd_pr__pfet_01v8_lvt_9UM225_0
timestamp 1663011646
transform 1 0 968 0 1 712
box -968 -712 968 745
<< end >>
