magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -971 -795 971 857
<< nmoslvt >>
rect -887 -769 -487 831
rect -429 -769 -29 831
rect 29 -769 429 831
rect 487 -769 887 831
<< ndiff >>
rect -945 796 -887 831
rect -945 762 -933 796
rect -899 762 -887 796
rect -945 728 -887 762
rect -945 694 -933 728
rect -899 694 -887 728
rect -945 660 -887 694
rect -945 626 -933 660
rect -899 626 -887 660
rect -945 592 -887 626
rect -945 558 -933 592
rect -899 558 -887 592
rect -945 524 -887 558
rect -945 490 -933 524
rect -899 490 -887 524
rect -945 456 -887 490
rect -945 422 -933 456
rect -899 422 -887 456
rect -945 388 -887 422
rect -945 354 -933 388
rect -899 354 -887 388
rect -945 320 -887 354
rect -945 286 -933 320
rect -899 286 -887 320
rect -945 252 -887 286
rect -945 218 -933 252
rect -899 218 -887 252
rect -945 184 -887 218
rect -945 150 -933 184
rect -899 150 -887 184
rect -945 116 -887 150
rect -945 82 -933 116
rect -899 82 -887 116
rect -945 48 -887 82
rect -945 14 -933 48
rect -899 14 -887 48
rect -945 -20 -887 14
rect -945 -54 -933 -20
rect -899 -54 -887 -20
rect -945 -88 -887 -54
rect -945 -122 -933 -88
rect -899 -122 -887 -88
rect -945 -156 -887 -122
rect -945 -190 -933 -156
rect -899 -190 -887 -156
rect -945 -224 -887 -190
rect -945 -258 -933 -224
rect -899 -258 -887 -224
rect -945 -292 -887 -258
rect -945 -326 -933 -292
rect -899 -326 -887 -292
rect -945 -360 -887 -326
rect -945 -394 -933 -360
rect -899 -394 -887 -360
rect -945 -428 -887 -394
rect -945 -462 -933 -428
rect -899 -462 -887 -428
rect -945 -496 -887 -462
rect -945 -530 -933 -496
rect -899 -530 -887 -496
rect -945 -564 -887 -530
rect -945 -598 -933 -564
rect -899 -598 -887 -564
rect -945 -632 -887 -598
rect -945 -666 -933 -632
rect -899 -666 -887 -632
rect -945 -700 -887 -666
rect -945 -734 -933 -700
rect -899 -734 -887 -700
rect -945 -769 -887 -734
rect -487 796 -429 831
rect -487 762 -475 796
rect -441 762 -429 796
rect -487 728 -429 762
rect -487 694 -475 728
rect -441 694 -429 728
rect -487 660 -429 694
rect -487 626 -475 660
rect -441 626 -429 660
rect -487 592 -429 626
rect -487 558 -475 592
rect -441 558 -429 592
rect -487 524 -429 558
rect -487 490 -475 524
rect -441 490 -429 524
rect -487 456 -429 490
rect -487 422 -475 456
rect -441 422 -429 456
rect -487 388 -429 422
rect -487 354 -475 388
rect -441 354 -429 388
rect -487 320 -429 354
rect -487 286 -475 320
rect -441 286 -429 320
rect -487 252 -429 286
rect -487 218 -475 252
rect -441 218 -429 252
rect -487 184 -429 218
rect -487 150 -475 184
rect -441 150 -429 184
rect -487 116 -429 150
rect -487 82 -475 116
rect -441 82 -429 116
rect -487 48 -429 82
rect -487 14 -475 48
rect -441 14 -429 48
rect -487 -20 -429 14
rect -487 -54 -475 -20
rect -441 -54 -429 -20
rect -487 -88 -429 -54
rect -487 -122 -475 -88
rect -441 -122 -429 -88
rect -487 -156 -429 -122
rect -487 -190 -475 -156
rect -441 -190 -429 -156
rect -487 -224 -429 -190
rect -487 -258 -475 -224
rect -441 -258 -429 -224
rect -487 -292 -429 -258
rect -487 -326 -475 -292
rect -441 -326 -429 -292
rect -487 -360 -429 -326
rect -487 -394 -475 -360
rect -441 -394 -429 -360
rect -487 -428 -429 -394
rect -487 -462 -475 -428
rect -441 -462 -429 -428
rect -487 -496 -429 -462
rect -487 -530 -475 -496
rect -441 -530 -429 -496
rect -487 -564 -429 -530
rect -487 -598 -475 -564
rect -441 -598 -429 -564
rect -487 -632 -429 -598
rect -487 -666 -475 -632
rect -441 -666 -429 -632
rect -487 -700 -429 -666
rect -487 -734 -475 -700
rect -441 -734 -429 -700
rect -487 -769 -429 -734
rect -29 796 29 831
rect -29 762 -17 796
rect 17 762 29 796
rect -29 728 29 762
rect -29 694 -17 728
rect 17 694 29 728
rect -29 660 29 694
rect -29 626 -17 660
rect 17 626 29 660
rect -29 592 29 626
rect -29 558 -17 592
rect 17 558 29 592
rect -29 524 29 558
rect -29 490 -17 524
rect 17 490 29 524
rect -29 456 29 490
rect -29 422 -17 456
rect 17 422 29 456
rect -29 388 29 422
rect -29 354 -17 388
rect 17 354 29 388
rect -29 320 29 354
rect -29 286 -17 320
rect 17 286 29 320
rect -29 252 29 286
rect -29 218 -17 252
rect 17 218 29 252
rect -29 184 29 218
rect -29 150 -17 184
rect 17 150 29 184
rect -29 116 29 150
rect -29 82 -17 116
rect 17 82 29 116
rect -29 48 29 82
rect -29 14 -17 48
rect 17 14 29 48
rect -29 -20 29 14
rect -29 -54 -17 -20
rect 17 -54 29 -20
rect -29 -88 29 -54
rect -29 -122 -17 -88
rect 17 -122 29 -88
rect -29 -156 29 -122
rect -29 -190 -17 -156
rect 17 -190 29 -156
rect -29 -224 29 -190
rect -29 -258 -17 -224
rect 17 -258 29 -224
rect -29 -292 29 -258
rect -29 -326 -17 -292
rect 17 -326 29 -292
rect -29 -360 29 -326
rect -29 -394 -17 -360
rect 17 -394 29 -360
rect -29 -428 29 -394
rect -29 -462 -17 -428
rect 17 -462 29 -428
rect -29 -496 29 -462
rect -29 -530 -17 -496
rect 17 -530 29 -496
rect -29 -564 29 -530
rect -29 -598 -17 -564
rect 17 -598 29 -564
rect -29 -632 29 -598
rect -29 -666 -17 -632
rect 17 -666 29 -632
rect -29 -700 29 -666
rect -29 -734 -17 -700
rect 17 -734 29 -700
rect -29 -769 29 -734
rect 429 796 487 831
rect 429 762 441 796
rect 475 762 487 796
rect 429 728 487 762
rect 429 694 441 728
rect 475 694 487 728
rect 429 660 487 694
rect 429 626 441 660
rect 475 626 487 660
rect 429 592 487 626
rect 429 558 441 592
rect 475 558 487 592
rect 429 524 487 558
rect 429 490 441 524
rect 475 490 487 524
rect 429 456 487 490
rect 429 422 441 456
rect 475 422 487 456
rect 429 388 487 422
rect 429 354 441 388
rect 475 354 487 388
rect 429 320 487 354
rect 429 286 441 320
rect 475 286 487 320
rect 429 252 487 286
rect 429 218 441 252
rect 475 218 487 252
rect 429 184 487 218
rect 429 150 441 184
rect 475 150 487 184
rect 429 116 487 150
rect 429 82 441 116
rect 475 82 487 116
rect 429 48 487 82
rect 429 14 441 48
rect 475 14 487 48
rect 429 -20 487 14
rect 429 -54 441 -20
rect 475 -54 487 -20
rect 429 -88 487 -54
rect 429 -122 441 -88
rect 475 -122 487 -88
rect 429 -156 487 -122
rect 429 -190 441 -156
rect 475 -190 487 -156
rect 429 -224 487 -190
rect 429 -258 441 -224
rect 475 -258 487 -224
rect 429 -292 487 -258
rect 429 -326 441 -292
rect 475 -326 487 -292
rect 429 -360 487 -326
rect 429 -394 441 -360
rect 475 -394 487 -360
rect 429 -428 487 -394
rect 429 -462 441 -428
rect 475 -462 487 -428
rect 429 -496 487 -462
rect 429 -530 441 -496
rect 475 -530 487 -496
rect 429 -564 487 -530
rect 429 -598 441 -564
rect 475 -598 487 -564
rect 429 -632 487 -598
rect 429 -666 441 -632
rect 475 -666 487 -632
rect 429 -700 487 -666
rect 429 -734 441 -700
rect 475 -734 487 -700
rect 429 -769 487 -734
rect 887 796 945 831
rect 887 762 899 796
rect 933 762 945 796
rect 887 728 945 762
rect 887 694 899 728
rect 933 694 945 728
rect 887 660 945 694
rect 887 626 899 660
rect 933 626 945 660
rect 887 592 945 626
rect 887 558 899 592
rect 933 558 945 592
rect 887 524 945 558
rect 887 490 899 524
rect 933 490 945 524
rect 887 456 945 490
rect 887 422 899 456
rect 933 422 945 456
rect 887 388 945 422
rect 887 354 899 388
rect 933 354 945 388
rect 887 320 945 354
rect 887 286 899 320
rect 933 286 945 320
rect 887 252 945 286
rect 887 218 899 252
rect 933 218 945 252
rect 887 184 945 218
rect 887 150 899 184
rect 933 150 945 184
rect 887 116 945 150
rect 887 82 899 116
rect 933 82 945 116
rect 887 48 945 82
rect 887 14 899 48
rect 933 14 945 48
rect 887 -20 945 14
rect 887 -54 899 -20
rect 933 -54 945 -20
rect 887 -88 945 -54
rect 887 -122 899 -88
rect 933 -122 945 -88
rect 887 -156 945 -122
rect 887 -190 899 -156
rect 933 -190 945 -156
rect 887 -224 945 -190
rect 887 -258 899 -224
rect 933 -258 945 -224
rect 887 -292 945 -258
rect 887 -326 899 -292
rect 933 -326 945 -292
rect 887 -360 945 -326
rect 887 -394 899 -360
rect 933 -394 945 -360
rect 887 -428 945 -394
rect 887 -462 899 -428
rect 933 -462 945 -428
rect 887 -496 945 -462
rect 887 -530 899 -496
rect 933 -530 945 -496
rect 887 -564 945 -530
rect 887 -598 899 -564
rect 933 -598 945 -564
rect 887 -632 945 -598
rect 887 -666 899 -632
rect 933 -666 945 -632
rect 887 -700 945 -666
rect 887 -734 899 -700
rect 933 -734 945 -700
rect 887 -769 945 -734
<< ndiffc >>
rect -933 762 -899 796
rect -933 694 -899 728
rect -933 626 -899 660
rect -933 558 -899 592
rect -933 490 -899 524
rect -933 422 -899 456
rect -933 354 -899 388
rect -933 286 -899 320
rect -933 218 -899 252
rect -933 150 -899 184
rect -933 82 -899 116
rect -933 14 -899 48
rect -933 -54 -899 -20
rect -933 -122 -899 -88
rect -933 -190 -899 -156
rect -933 -258 -899 -224
rect -933 -326 -899 -292
rect -933 -394 -899 -360
rect -933 -462 -899 -428
rect -933 -530 -899 -496
rect -933 -598 -899 -564
rect -933 -666 -899 -632
rect -933 -734 -899 -700
rect -475 762 -441 796
rect -475 694 -441 728
rect -475 626 -441 660
rect -475 558 -441 592
rect -475 490 -441 524
rect -475 422 -441 456
rect -475 354 -441 388
rect -475 286 -441 320
rect -475 218 -441 252
rect -475 150 -441 184
rect -475 82 -441 116
rect -475 14 -441 48
rect -475 -54 -441 -20
rect -475 -122 -441 -88
rect -475 -190 -441 -156
rect -475 -258 -441 -224
rect -475 -326 -441 -292
rect -475 -394 -441 -360
rect -475 -462 -441 -428
rect -475 -530 -441 -496
rect -475 -598 -441 -564
rect -475 -666 -441 -632
rect -475 -734 -441 -700
rect -17 762 17 796
rect -17 694 17 728
rect -17 626 17 660
rect -17 558 17 592
rect -17 490 17 524
rect -17 422 17 456
rect -17 354 17 388
rect -17 286 17 320
rect -17 218 17 252
rect -17 150 17 184
rect -17 82 17 116
rect -17 14 17 48
rect -17 -54 17 -20
rect -17 -122 17 -88
rect -17 -190 17 -156
rect -17 -258 17 -224
rect -17 -326 17 -292
rect -17 -394 17 -360
rect -17 -462 17 -428
rect -17 -530 17 -496
rect -17 -598 17 -564
rect -17 -666 17 -632
rect -17 -734 17 -700
rect 441 762 475 796
rect 441 694 475 728
rect 441 626 475 660
rect 441 558 475 592
rect 441 490 475 524
rect 441 422 475 456
rect 441 354 475 388
rect 441 286 475 320
rect 441 218 475 252
rect 441 150 475 184
rect 441 82 475 116
rect 441 14 475 48
rect 441 -54 475 -20
rect 441 -122 475 -88
rect 441 -190 475 -156
rect 441 -258 475 -224
rect 441 -326 475 -292
rect 441 -394 475 -360
rect 441 -462 475 -428
rect 441 -530 475 -496
rect 441 -598 475 -564
rect 441 -666 475 -632
rect 441 -734 475 -700
rect 899 762 933 796
rect 899 694 933 728
rect 899 626 933 660
rect 899 558 933 592
rect 899 490 933 524
rect 899 422 933 456
rect 899 354 933 388
rect 899 286 933 320
rect 899 218 933 252
rect 899 150 933 184
rect 899 82 933 116
rect 899 14 933 48
rect 899 -54 933 -20
rect 899 -122 933 -88
rect 899 -190 933 -156
rect 899 -258 933 -224
rect 899 -326 933 -292
rect 899 -394 933 -360
rect 899 -462 933 -428
rect 899 -530 933 -496
rect 899 -598 933 -564
rect 899 -666 933 -632
rect 899 -734 933 -700
<< poly >>
rect -887 831 -487 857
rect -429 831 -29 857
rect 29 831 429 857
rect 487 831 887 857
rect -887 -807 -487 -769
rect -887 -841 -840 -807
rect -806 -841 -772 -807
rect -738 -841 -704 -807
rect -670 -841 -636 -807
rect -602 -841 -568 -807
rect -534 -841 -487 -807
rect -887 -857 -487 -841
rect -429 -807 -29 -769
rect -429 -841 -382 -807
rect -348 -841 -314 -807
rect -280 -841 -246 -807
rect -212 -841 -178 -807
rect -144 -841 -110 -807
rect -76 -841 -29 -807
rect -429 -857 -29 -841
rect 29 -807 429 -769
rect 29 -841 76 -807
rect 110 -841 144 -807
rect 178 -841 212 -807
rect 246 -841 280 -807
rect 314 -841 348 -807
rect 382 -841 429 -807
rect 29 -857 429 -841
rect 487 -807 887 -769
rect 487 -841 534 -807
rect 568 -841 602 -807
rect 636 -841 670 -807
rect 704 -841 738 -807
rect 772 -841 806 -807
rect 840 -841 887 -807
rect 487 -857 887 -841
<< polycont >>
rect -840 -841 -806 -807
rect -772 -841 -738 -807
rect -704 -841 -670 -807
rect -636 -841 -602 -807
rect -568 -841 -534 -807
rect -382 -841 -348 -807
rect -314 -841 -280 -807
rect -246 -841 -212 -807
rect -178 -841 -144 -807
rect -110 -841 -76 -807
rect 76 -841 110 -807
rect 144 -841 178 -807
rect 212 -841 246 -807
rect 280 -841 314 -807
rect 348 -841 382 -807
rect 534 -841 568 -807
rect 602 -841 636 -807
rect 670 -841 704 -807
rect 738 -841 772 -807
rect 806 -841 840 -807
<< locali >>
rect -933 804 -899 835
rect -933 732 -899 762
rect -933 660 -899 694
rect -933 592 -899 626
rect -933 524 -899 554
rect -933 456 -899 482
rect -933 388 -899 410
rect -933 320 -899 338
rect -933 252 -899 266
rect -933 184 -899 194
rect -933 116 -899 122
rect -933 48 -899 50
rect -933 12 -899 14
rect -933 -60 -899 -54
rect -933 -132 -899 -122
rect -933 -204 -899 -190
rect -933 -276 -899 -258
rect -933 -348 -899 -326
rect -933 -420 -899 -394
rect -933 -492 -899 -462
rect -933 -564 -899 -530
rect -933 -632 -899 -598
rect -933 -700 -899 -670
rect -933 -773 -899 -742
rect -475 804 -441 835
rect -475 732 -441 762
rect -475 660 -441 694
rect -475 592 -441 626
rect -475 524 -441 554
rect -475 456 -441 482
rect -475 388 -441 410
rect -475 320 -441 338
rect -475 252 -441 266
rect -475 184 -441 194
rect -475 116 -441 122
rect -475 48 -441 50
rect -475 12 -441 14
rect -475 -60 -441 -54
rect -475 -132 -441 -122
rect -475 -204 -441 -190
rect -475 -276 -441 -258
rect -475 -348 -441 -326
rect -475 -420 -441 -394
rect -475 -492 -441 -462
rect -475 -564 -441 -530
rect -475 -632 -441 -598
rect -475 -700 -441 -670
rect -475 -773 -441 -742
rect -17 804 17 835
rect -17 732 17 762
rect -17 660 17 694
rect -17 592 17 626
rect -17 524 17 554
rect -17 456 17 482
rect -17 388 17 410
rect -17 320 17 338
rect -17 252 17 266
rect -17 184 17 194
rect -17 116 17 122
rect -17 48 17 50
rect -17 12 17 14
rect -17 -60 17 -54
rect -17 -132 17 -122
rect -17 -204 17 -190
rect -17 -276 17 -258
rect -17 -348 17 -326
rect -17 -420 17 -394
rect -17 -492 17 -462
rect -17 -564 17 -530
rect -17 -632 17 -598
rect -17 -700 17 -670
rect -17 -773 17 -742
rect 441 804 475 835
rect 441 732 475 762
rect 441 660 475 694
rect 441 592 475 626
rect 441 524 475 554
rect 441 456 475 482
rect 441 388 475 410
rect 441 320 475 338
rect 441 252 475 266
rect 441 184 475 194
rect 441 116 475 122
rect 441 48 475 50
rect 441 12 475 14
rect 441 -60 475 -54
rect 441 -132 475 -122
rect 441 -204 475 -190
rect 441 -276 475 -258
rect 441 -348 475 -326
rect 441 -420 475 -394
rect 441 -492 475 -462
rect 441 -564 475 -530
rect 441 -632 475 -598
rect 441 -700 475 -670
rect 441 -773 475 -742
rect 899 804 933 835
rect 899 732 933 762
rect 899 660 933 694
rect 899 592 933 626
rect 899 524 933 554
rect 899 456 933 482
rect 899 388 933 410
rect 899 320 933 338
rect 899 252 933 266
rect 899 184 933 194
rect 899 116 933 122
rect 899 48 933 50
rect 899 12 933 14
rect 899 -60 933 -54
rect 899 -132 933 -122
rect 899 -204 933 -190
rect 899 -276 933 -258
rect 899 -348 933 -326
rect 899 -420 933 -394
rect 899 -492 933 -462
rect 899 -564 933 -530
rect 899 -632 933 -598
rect 899 -700 933 -670
rect 899 -773 933 -742
rect -887 -841 -848 -807
rect -806 -841 -776 -807
rect -738 -841 -704 -807
rect -670 -841 -636 -807
rect -598 -841 -568 -807
rect -526 -841 -487 -807
rect -429 -841 -390 -807
rect -348 -841 -318 -807
rect -280 -841 -246 -807
rect -212 -841 -178 -807
rect -140 -841 -110 -807
rect -68 -841 -29 -807
rect 29 -841 68 -807
rect 110 -841 140 -807
rect 178 -841 212 -807
rect 246 -841 280 -807
rect 318 -841 348 -807
rect 390 -841 429 -807
rect 487 -841 526 -807
rect 568 -841 598 -807
rect 636 -841 670 -807
rect 704 -841 738 -807
rect 776 -841 806 -807
rect 848 -841 887 -807
<< viali >>
rect -933 796 -899 804
rect -933 770 -899 796
rect -933 728 -899 732
rect -933 698 -899 728
rect -933 626 -899 660
rect -933 558 -899 588
rect -933 554 -899 558
rect -933 490 -899 516
rect -933 482 -899 490
rect -933 422 -899 444
rect -933 410 -899 422
rect -933 354 -899 372
rect -933 338 -899 354
rect -933 286 -899 300
rect -933 266 -899 286
rect -933 218 -899 228
rect -933 194 -899 218
rect -933 150 -899 156
rect -933 122 -899 150
rect -933 82 -899 84
rect -933 50 -899 82
rect -933 -20 -899 12
rect -933 -22 -899 -20
rect -933 -88 -899 -60
rect -933 -94 -899 -88
rect -933 -156 -899 -132
rect -933 -166 -899 -156
rect -933 -224 -899 -204
rect -933 -238 -899 -224
rect -933 -292 -899 -276
rect -933 -310 -899 -292
rect -933 -360 -899 -348
rect -933 -382 -899 -360
rect -933 -428 -899 -420
rect -933 -454 -899 -428
rect -933 -496 -899 -492
rect -933 -526 -899 -496
rect -933 -598 -899 -564
rect -933 -666 -899 -636
rect -933 -670 -899 -666
rect -933 -734 -899 -708
rect -933 -742 -899 -734
rect -475 796 -441 804
rect -475 770 -441 796
rect -475 728 -441 732
rect -475 698 -441 728
rect -475 626 -441 660
rect -475 558 -441 588
rect -475 554 -441 558
rect -475 490 -441 516
rect -475 482 -441 490
rect -475 422 -441 444
rect -475 410 -441 422
rect -475 354 -441 372
rect -475 338 -441 354
rect -475 286 -441 300
rect -475 266 -441 286
rect -475 218 -441 228
rect -475 194 -441 218
rect -475 150 -441 156
rect -475 122 -441 150
rect -475 82 -441 84
rect -475 50 -441 82
rect -475 -20 -441 12
rect -475 -22 -441 -20
rect -475 -88 -441 -60
rect -475 -94 -441 -88
rect -475 -156 -441 -132
rect -475 -166 -441 -156
rect -475 -224 -441 -204
rect -475 -238 -441 -224
rect -475 -292 -441 -276
rect -475 -310 -441 -292
rect -475 -360 -441 -348
rect -475 -382 -441 -360
rect -475 -428 -441 -420
rect -475 -454 -441 -428
rect -475 -496 -441 -492
rect -475 -526 -441 -496
rect -475 -598 -441 -564
rect -475 -666 -441 -636
rect -475 -670 -441 -666
rect -475 -734 -441 -708
rect -475 -742 -441 -734
rect -17 796 17 804
rect -17 770 17 796
rect -17 728 17 732
rect -17 698 17 728
rect -17 626 17 660
rect -17 558 17 588
rect -17 554 17 558
rect -17 490 17 516
rect -17 482 17 490
rect -17 422 17 444
rect -17 410 17 422
rect -17 354 17 372
rect -17 338 17 354
rect -17 286 17 300
rect -17 266 17 286
rect -17 218 17 228
rect -17 194 17 218
rect -17 150 17 156
rect -17 122 17 150
rect -17 82 17 84
rect -17 50 17 82
rect -17 -20 17 12
rect -17 -22 17 -20
rect -17 -88 17 -60
rect -17 -94 17 -88
rect -17 -156 17 -132
rect -17 -166 17 -156
rect -17 -224 17 -204
rect -17 -238 17 -224
rect -17 -292 17 -276
rect -17 -310 17 -292
rect -17 -360 17 -348
rect -17 -382 17 -360
rect -17 -428 17 -420
rect -17 -454 17 -428
rect -17 -496 17 -492
rect -17 -526 17 -496
rect -17 -598 17 -564
rect -17 -666 17 -636
rect -17 -670 17 -666
rect -17 -734 17 -708
rect -17 -742 17 -734
rect 441 796 475 804
rect 441 770 475 796
rect 441 728 475 732
rect 441 698 475 728
rect 441 626 475 660
rect 441 558 475 588
rect 441 554 475 558
rect 441 490 475 516
rect 441 482 475 490
rect 441 422 475 444
rect 441 410 475 422
rect 441 354 475 372
rect 441 338 475 354
rect 441 286 475 300
rect 441 266 475 286
rect 441 218 475 228
rect 441 194 475 218
rect 441 150 475 156
rect 441 122 475 150
rect 441 82 475 84
rect 441 50 475 82
rect 441 -20 475 12
rect 441 -22 475 -20
rect 441 -88 475 -60
rect 441 -94 475 -88
rect 441 -156 475 -132
rect 441 -166 475 -156
rect 441 -224 475 -204
rect 441 -238 475 -224
rect 441 -292 475 -276
rect 441 -310 475 -292
rect 441 -360 475 -348
rect 441 -382 475 -360
rect 441 -428 475 -420
rect 441 -454 475 -428
rect 441 -496 475 -492
rect 441 -526 475 -496
rect 441 -598 475 -564
rect 441 -666 475 -636
rect 441 -670 475 -666
rect 441 -734 475 -708
rect 441 -742 475 -734
rect 899 796 933 804
rect 899 770 933 796
rect 899 728 933 732
rect 899 698 933 728
rect 899 626 933 660
rect 899 558 933 588
rect 899 554 933 558
rect 899 490 933 516
rect 899 482 933 490
rect 899 422 933 444
rect 899 410 933 422
rect 899 354 933 372
rect 899 338 933 354
rect 899 286 933 300
rect 899 266 933 286
rect 899 218 933 228
rect 899 194 933 218
rect 899 150 933 156
rect 899 122 933 150
rect 899 82 933 84
rect 899 50 933 82
rect 899 -20 933 12
rect 899 -22 933 -20
rect 899 -88 933 -60
rect 899 -94 933 -88
rect 899 -156 933 -132
rect 899 -166 933 -156
rect 899 -224 933 -204
rect 899 -238 933 -224
rect 899 -292 933 -276
rect 899 -310 933 -292
rect 899 -360 933 -348
rect 899 -382 933 -360
rect 899 -428 933 -420
rect 899 -454 933 -428
rect 899 -496 933 -492
rect 899 -526 933 -496
rect 899 -598 933 -564
rect 899 -666 933 -636
rect 899 -670 933 -666
rect 899 -734 933 -708
rect 899 -742 933 -734
rect -848 -841 -840 -807
rect -840 -841 -814 -807
rect -776 -841 -772 -807
rect -772 -841 -742 -807
rect -704 -841 -670 -807
rect -632 -841 -602 -807
rect -602 -841 -598 -807
rect -560 -841 -534 -807
rect -534 -841 -526 -807
rect -390 -841 -382 -807
rect -382 -841 -356 -807
rect -318 -841 -314 -807
rect -314 -841 -284 -807
rect -246 -841 -212 -807
rect -174 -841 -144 -807
rect -144 -841 -140 -807
rect -102 -841 -76 -807
rect -76 -841 -68 -807
rect 68 -841 76 -807
rect 76 -841 102 -807
rect 140 -841 144 -807
rect 144 -841 174 -807
rect 212 -841 246 -807
rect 284 -841 314 -807
rect 314 -841 318 -807
rect 356 -841 382 -807
rect 382 -841 390 -807
rect 526 -841 534 -807
rect 534 -841 560 -807
rect 598 -841 602 -807
rect 602 -841 632 -807
rect 670 -841 704 -807
rect 742 -841 772 -807
rect 772 -841 776 -807
rect 814 -841 840 -807
rect 840 -841 848 -807
<< metal1 >>
rect -939 804 -893 831
rect -939 770 -933 804
rect -899 770 -893 804
rect -939 732 -893 770
rect -939 698 -933 732
rect -899 698 -893 732
rect -939 660 -893 698
rect -939 626 -933 660
rect -899 626 -893 660
rect -939 588 -893 626
rect -939 554 -933 588
rect -899 554 -893 588
rect -939 516 -893 554
rect -939 482 -933 516
rect -899 482 -893 516
rect -939 444 -893 482
rect -939 410 -933 444
rect -899 410 -893 444
rect -939 372 -893 410
rect -939 338 -933 372
rect -899 338 -893 372
rect -939 300 -893 338
rect -939 266 -933 300
rect -899 266 -893 300
rect -939 228 -893 266
rect -939 194 -933 228
rect -899 194 -893 228
rect -939 156 -893 194
rect -939 122 -933 156
rect -899 122 -893 156
rect -939 84 -893 122
rect -939 50 -933 84
rect -899 50 -893 84
rect -939 12 -893 50
rect -939 -22 -933 12
rect -899 -22 -893 12
rect -939 -60 -893 -22
rect -939 -94 -933 -60
rect -899 -94 -893 -60
rect -939 -132 -893 -94
rect -939 -166 -933 -132
rect -899 -166 -893 -132
rect -939 -204 -893 -166
rect -939 -238 -933 -204
rect -899 -238 -893 -204
rect -939 -276 -893 -238
rect -939 -310 -933 -276
rect -899 -310 -893 -276
rect -939 -348 -893 -310
rect -939 -382 -933 -348
rect -899 -382 -893 -348
rect -939 -420 -893 -382
rect -939 -454 -933 -420
rect -899 -454 -893 -420
rect -939 -492 -893 -454
rect -939 -526 -933 -492
rect -899 -526 -893 -492
rect -939 -564 -893 -526
rect -939 -598 -933 -564
rect -899 -598 -893 -564
rect -939 -636 -893 -598
rect -939 -670 -933 -636
rect -899 -670 -893 -636
rect -939 -708 -893 -670
rect -939 -742 -933 -708
rect -899 -742 -893 -708
rect -939 -769 -893 -742
rect -481 804 -435 831
rect -481 770 -475 804
rect -441 770 -435 804
rect -481 732 -435 770
rect -481 698 -475 732
rect -441 698 -435 732
rect -481 660 -435 698
rect -481 626 -475 660
rect -441 626 -435 660
rect -481 588 -435 626
rect -481 554 -475 588
rect -441 554 -435 588
rect -481 516 -435 554
rect -481 482 -475 516
rect -441 482 -435 516
rect -481 444 -435 482
rect -481 410 -475 444
rect -441 410 -435 444
rect -481 372 -435 410
rect -481 338 -475 372
rect -441 338 -435 372
rect -481 300 -435 338
rect -481 266 -475 300
rect -441 266 -435 300
rect -481 228 -435 266
rect -481 194 -475 228
rect -441 194 -435 228
rect -481 156 -435 194
rect -481 122 -475 156
rect -441 122 -435 156
rect -481 84 -435 122
rect -481 50 -475 84
rect -441 50 -435 84
rect -481 12 -435 50
rect -481 -22 -475 12
rect -441 -22 -435 12
rect -481 -60 -435 -22
rect -481 -94 -475 -60
rect -441 -94 -435 -60
rect -481 -132 -435 -94
rect -481 -166 -475 -132
rect -441 -166 -435 -132
rect -481 -204 -435 -166
rect -481 -238 -475 -204
rect -441 -238 -435 -204
rect -481 -276 -435 -238
rect -481 -310 -475 -276
rect -441 -310 -435 -276
rect -481 -348 -435 -310
rect -481 -382 -475 -348
rect -441 -382 -435 -348
rect -481 -420 -435 -382
rect -481 -454 -475 -420
rect -441 -454 -435 -420
rect -481 -492 -435 -454
rect -481 -526 -475 -492
rect -441 -526 -435 -492
rect -481 -564 -435 -526
rect -481 -598 -475 -564
rect -441 -598 -435 -564
rect -481 -636 -435 -598
rect -481 -670 -475 -636
rect -441 -670 -435 -636
rect -481 -708 -435 -670
rect -481 -742 -475 -708
rect -441 -742 -435 -708
rect -481 -769 -435 -742
rect -23 804 23 831
rect -23 770 -17 804
rect 17 770 23 804
rect -23 732 23 770
rect -23 698 -17 732
rect 17 698 23 732
rect -23 660 23 698
rect -23 626 -17 660
rect 17 626 23 660
rect -23 588 23 626
rect -23 554 -17 588
rect 17 554 23 588
rect -23 516 23 554
rect -23 482 -17 516
rect 17 482 23 516
rect -23 444 23 482
rect -23 410 -17 444
rect 17 410 23 444
rect -23 372 23 410
rect -23 338 -17 372
rect 17 338 23 372
rect -23 300 23 338
rect -23 266 -17 300
rect 17 266 23 300
rect -23 228 23 266
rect -23 194 -17 228
rect 17 194 23 228
rect -23 156 23 194
rect -23 122 -17 156
rect 17 122 23 156
rect -23 84 23 122
rect -23 50 -17 84
rect 17 50 23 84
rect -23 12 23 50
rect -23 -22 -17 12
rect 17 -22 23 12
rect -23 -60 23 -22
rect -23 -94 -17 -60
rect 17 -94 23 -60
rect -23 -132 23 -94
rect -23 -166 -17 -132
rect 17 -166 23 -132
rect -23 -204 23 -166
rect -23 -238 -17 -204
rect 17 -238 23 -204
rect -23 -276 23 -238
rect -23 -310 -17 -276
rect 17 -310 23 -276
rect -23 -348 23 -310
rect -23 -382 -17 -348
rect 17 -382 23 -348
rect -23 -420 23 -382
rect -23 -454 -17 -420
rect 17 -454 23 -420
rect -23 -492 23 -454
rect -23 -526 -17 -492
rect 17 -526 23 -492
rect -23 -564 23 -526
rect -23 -598 -17 -564
rect 17 -598 23 -564
rect -23 -636 23 -598
rect -23 -670 -17 -636
rect 17 -670 23 -636
rect -23 -708 23 -670
rect -23 -742 -17 -708
rect 17 -742 23 -708
rect -23 -769 23 -742
rect 435 804 481 831
rect 435 770 441 804
rect 475 770 481 804
rect 435 732 481 770
rect 435 698 441 732
rect 475 698 481 732
rect 435 660 481 698
rect 435 626 441 660
rect 475 626 481 660
rect 435 588 481 626
rect 435 554 441 588
rect 475 554 481 588
rect 435 516 481 554
rect 435 482 441 516
rect 475 482 481 516
rect 435 444 481 482
rect 435 410 441 444
rect 475 410 481 444
rect 435 372 481 410
rect 435 338 441 372
rect 475 338 481 372
rect 435 300 481 338
rect 435 266 441 300
rect 475 266 481 300
rect 435 228 481 266
rect 435 194 441 228
rect 475 194 481 228
rect 435 156 481 194
rect 435 122 441 156
rect 475 122 481 156
rect 435 84 481 122
rect 435 50 441 84
rect 475 50 481 84
rect 435 12 481 50
rect 435 -22 441 12
rect 475 -22 481 12
rect 435 -60 481 -22
rect 435 -94 441 -60
rect 475 -94 481 -60
rect 435 -132 481 -94
rect 435 -166 441 -132
rect 475 -166 481 -132
rect 435 -204 481 -166
rect 435 -238 441 -204
rect 475 -238 481 -204
rect 435 -276 481 -238
rect 435 -310 441 -276
rect 475 -310 481 -276
rect 435 -348 481 -310
rect 435 -382 441 -348
rect 475 -382 481 -348
rect 435 -420 481 -382
rect 435 -454 441 -420
rect 475 -454 481 -420
rect 435 -492 481 -454
rect 435 -526 441 -492
rect 475 -526 481 -492
rect 435 -564 481 -526
rect 435 -598 441 -564
rect 475 -598 481 -564
rect 435 -636 481 -598
rect 435 -670 441 -636
rect 475 -670 481 -636
rect 435 -708 481 -670
rect 435 -742 441 -708
rect 475 -742 481 -708
rect 435 -769 481 -742
rect 893 804 939 831
rect 893 770 899 804
rect 933 770 939 804
rect 893 732 939 770
rect 893 698 899 732
rect 933 698 939 732
rect 893 660 939 698
rect 893 626 899 660
rect 933 626 939 660
rect 893 588 939 626
rect 893 554 899 588
rect 933 554 939 588
rect 893 516 939 554
rect 893 482 899 516
rect 933 482 939 516
rect 893 444 939 482
rect 893 410 899 444
rect 933 410 939 444
rect 893 372 939 410
rect 893 338 899 372
rect 933 338 939 372
rect 893 300 939 338
rect 893 266 899 300
rect 933 266 939 300
rect 893 228 939 266
rect 893 194 899 228
rect 933 194 939 228
rect 893 156 939 194
rect 893 122 899 156
rect 933 122 939 156
rect 893 84 939 122
rect 893 50 899 84
rect 933 50 939 84
rect 893 12 939 50
rect 893 -22 899 12
rect 933 -22 939 12
rect 893 -60 939 -22
rect 893 -94 899 -60
rect 933 -94 939 -60
rect 893 -132 939 -94
rect 893 -166 899 -132
rect 933 -166 939 -132
rect 893 -204 939 -166
rect 893 -238 899 -204
rect 933 -238 939 -204
rect 893 -276 939 -238
rect 893 -310 899 -276
rect 933 -310 939 -276
rect 893 -348 939 -310
rect 893 -382 899 -348
rect 933 -382 939 -348
rect 893 -420 939 -382
rect 893 -454 899 -420
rect 933 -454 939 -420
rect 893 -492 939 -454
rect 893 -526 899 -492
rect 933 -526 939 -492
rect 893 -564 939 -526
rect 893 -598 899 -564
rect 933 -598 939 -564
rect 893 -636 939 -598
rect 893 -670 899 -636
rect 933 -670 939 -636
rect 893 -708 939 -670
rect 893 -742 899 -708
rect 933 -742 939 -708
rect 893 -769 939 -742
rect -883 -807 -491 -801
rect -883 -841 -848 -807
rect -814 -841 -776 -807
rect -742 -841 -704 -807
rect -670 -841 -632 -807
rect -598 -841 -560 -807
rect -526 -841 -491 -807
rect -883 -847 -491 -841
rect -425 -807 -33 -801
rect -425 -841 -390 -807
rect -356 -841 -318 -807
rect -284 -841 -246 -807
rect -212 -841 -174 -807
rect -140 -841 -102 -807
rect -68 -841 -33 -807
rect -425 -847 -33 -841
rect 33 -807 425 -801
rect 33 -841 68 -807
rect 102 -841 140 -807
rect 174 -841 212 -807
rect 246 -841 284 -807
rect 318 -841 356 -807
rect 390 -841 425 -807
rect 33 -847 425 -841
rect 491 -807 883 -801
rect 491 -841 526 -807
rect 560 -841 598 -807
rect 632 -841 670 -807
rect 704 -841 742 -807
rect 776 -841 814 -807
rect 848 -841 883 -807
rect 491 -847 883 -841
<< end >>
