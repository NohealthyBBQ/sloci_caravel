magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< nwell >>
rect -246 -584 246 584
<< pmos >>
rect -50 -364 50 436
<< pdiff >>
rect -108 393 -50 436
rect -108 359 -96 393
rect -62 359 -50 393
rect -108 325 -50 359
rect -108 291 -96 325
rect -62 291 -50 325
rect -108 257 -50 291
rect -108 223 -96 257
rect -62 223 -50 257
rect -108 189 -50 223
rect -108 155 -96 189
rect -62 155 -50 189
rect -108 121 -50 155
rect -108 87 -96 121
rect -62 87 -50 121
rect -108 53 -50 87
rect -108 19 -96 53
rect -62 19 -50 53
rect -108 -15 -50 19
rect -108 -49 -96 -15
rect -62 -49 -50 -15
rect -108 -83 -50 -49
rect -108 -117 -96 -83
rect -62 -117 -50 -83
rect -108 -151 -50 -117
rect -108 -185 -96 -151
rect -62 -185 -50 -151
rect -108 -219 -50 -185
rect -108 -253 -96 -219
rect -62 -253 -50 -219
rect -108 -287 -50 -253
rect -108 -321 -96 -287
rect -62 -321 -50 -287
rect -108 -364 -50 -321
rect 50 393 108 436
rect 50 359 62 393
rect 96 359 108 393
rect 50 325 108 359
rect 50 291 62 325
rect 96 291 108 325
rect 50 257 108 291
rect 50 223 62 257
rect 96 223 108 257
rect 50 189 108 223
rect 50 155 62 189
rect 96 155 108 189
rect 50 121 108 155
rect 50 87 62 121
rect 96 87 108 121
rect 50 53 108 87
rect 50 19 62 53
rect 96 19 108 53
rect 50 -15 108 19
rect 50 -49 62 -15
rect 96 -49 108 -15
rect 50 -83 108 -49
rect 50 -117 62 -83
rect 96 -117 108 -83
rect 50 -151 108 -117
rect 50 -185 62 -151
rect 96 -185 108 -151
rect 50 -219 108 -185
rect 50 -253 62 -219
rect 96 -253 108 -219
rect 50 -287 108 -253
rect 50 -321 62 -287
rect 96 -321 108 -287
rect 50 -364 108 -321
<< pdiffc >>
rect -96 359 -62 393
rect -96 291 -62 325
rect -96 223 -62 257
rect -96 155 -62 189
rect -96 87 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -15
rect -96 -117 -62 -83
rect -96 -185 -62 -151
rect -96 -253 -62 -219
rect -96 -321 -62 -287
rect 62 359 96 393
rect 62 291 96 325
rect 62 223 96 257
rect 62 155 96 189
rect 62 87 96 121
rect 62 19 96 53
rect 62 -49 96 -15
rect 62 -117 96 -83
rect 62 -185 96 -151
rect 62 -253 96 -219
rect 62 -321 96 -287
<< nsubdiff >>
rect -210 514 -85 548
rect -51 514 -17 548
rect 17 514 51 548
rect 85 514 210 548
rect -210 -514 -176 514
rect 176 -514 210 514
rect -210 -548 -85 -514
rect -51 -548 -17 -514
rect 17 -548 51 -514
rect 85 -548 210 -514
<< nsubdiffcont >>
rect -85 514 -51 548
rect -17 514 17 548
rect 51 514 85 548
rect -85 -548 -51 -514
rect -17 -548 17 -514
rect 51 -548 85 -514
<< poly >>
rect -50 436 50 462
rect -50 -411 50 -364
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect -50 -461 50 -445
<< polycont >>
rect -17 -445 17 -411
<< locali >>
rect -210 514 -85 548
rect -51 514 -17 548
rect 17 514 51 548
rect 85 514 210 548
rect -210 -514 -176 514
rect -96 413 -62 440
rect -96 341 -62 359
rect -96 269 -62 291
rect -96 197 -62 223
rect -96 125 -62 155
rect -96 53 -62 87
rect -96 -15 -62 19
rect -96 -83 -62 -53
rect -96 -151 -62 -125
rect -96 -219 -62 -197
rect -96 -287 -62 -269
rect -96 -368 -62 -341
rect 62 413 96 440
rect 62 341 96 359
rect 62 269 96 291
rect 62 197 96 223
rect 62 125 96 155
rect 62 53 96 87
rect 62 -15 96 19
rect 62 -83 96 -53
rect 62 -151 96 -125
rect 62 -219 96 -197
rect 62 -287 96 -269
rect 62 -368 96 -341
rect -50 -445 -17 -411
rect 17 -445 50 -411
rect 176 -514 210 514
rect -210 -548 -85 -514
rect -51 -548 -17 -514
rect 17 -548 51 -514
rect 85 -548 210 -514
<< viali >>
rect -96 393 -62 413
rect -96 379 -62 393
rect -96 325 -62 341
rect -96 307 -62 325
rect -96 257 -62 269
rect -96 235 -62 257
rect -96 189 -62 197
rect -96 163 -62 189
rect -96 121 -62 125
rect -96 91 -62 121
rect -96 19 -62 53
rect -96 -49 -62 -19
rect -96 -53 -62 -49
rect -96 -117 -62 -91
rect -96 -125 -62 -117
rect -96 -185 -62 -163
rect -96 -197 -62 -185
rect -96 -253 -62 -235
rect -96 -269 -62 -253
rect -96 -321 -62 -307
rect -96 -341 -62 -321
rect 62 393 96 413
rect 62 379 96 393
rect 62 325 96 341
rect 62 307 96 325
rect 62 257 96 269
rect 62 235 96 257
rect 62 189 96 197
rect 62 163 96 189
rect 62 121 96 125
rect 62 91 96 121
rect 62 19 96 53
rect 62 -49 96 -19
rect 62 -53 96 -49
rect 62 -117 96 -91
rect 62 -125 96 -117
rect 62 -185 96 -163
rect 62 -197 96 -185
rect 62 -253 96 -235
rect 62 -269 96 -253
rect 62 -321 96 -307
rect 62 -341 96 -321
rect -17 -445 17 -411
<< metal1 >>
rect -102 413 -56 436
rect -102 379 -96 413
rect -62 379 -56 413
rect -102 341 -56 379
rect -102 307 -96 341
rect -62 307 -56 341
rect -102 269 -56 307
rect -102 235 -96 269
rect -62 235 -56 269
rect -102 197 -56 235
rect -102 163 -96 197
rect -62 163 -56 197
rect -102 125 -56 163
rect -102 91 -96 125
rect -62 91 -56 125
rect -102 53 -56 91
rect -102 19 -96 53
rect -62 19 -56 53
rect -102 -19 -56 19
rect -102 -53 -96 -19
rect -62 -53 -56 -19
rect -102 -91 -56 -53
rect -102 -125 -96 -91
rect -62 -125 -56 -91
rect -102 -163 -56 -125
rect -102 -197 -96 -163
rect -62 -197 -56 -163
rect -102 -235 -56 -197
rect -102 -269 -96 -235
rect -62 -269 -56 -235
rect -102 -307 -56 -269
rect -102 -341 -96 -307
rect -62 -341 -56 -307
rect -102 -364 -56 -341
rect 56 413 102 436
rect 56 379 62 413
rect 96 379 102 413
rect 56 341 102 379
rect 56 307 62 341
rect 96 307 102 341
rect 56 269 102 307
rect 56 235 62 269
rect 96 235 102 269
rect 56 197 102 235
rect 56 163 62 197
rect 96 163 102 197
rect 56 125 102 163
rect 56 91 62 125
rect 96 91 102 125
rect 56 53 102 91
rect 56 19 62 53
rect 96 19 102 53
rect 56 -19 102 19
rect 56 -53 62 -19
rect 96 -53 102 -19
rect 56 -91 102 -53
rect 56 -125 62 -91
rect 96 -125 102 -91
rect 56 -163 102 -125
rect 56 -197 62 -163
rect 96 -197 102 -163
rect 56 -235 102 -197
rect 56 -269 62 -235
rect 96 -269 102 -235
rect 56 -307 102 -269
rect 56 -341 62 -307
rect 96 -341 102 -307
rect 56 -364 102 -341
rect -46 -411 46 -405
rect -46 -445 -17 -411
rect 17 -445 46 -411
rect -46 -451 46 -445
<< properties >>
string FIXED_BBOX -193 -531 193 531
<< end >>
