magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< locali >>
rect 6430 9730 6730 9770
rect 6430 8350 6730 8390
<< metal1 >>
rect 5770 9801 6340 9830
rect 5770 9429 5800 9801
rect 6300 9429 6340 9801
rect 5770 9400 6340 9429
rect 6780 8400 6840 9670
rect 6870 9666 7070 9670
rect 6870 9614 7004 9666
rect 7056 9614 7070 9666
rect 6870 9610 7070 9614
rect 6990 9600 7070 9610
rect 6870 9566 7070 9570
rect 6870 9514 6884 9566
rect 6936 9520 7070 9566
rect 6936 9514 6950 9520
rect 6870 9500 6950 9514
rect 6990 9476 7070 9480
rect 6990 9470 7004 9476
rect 6870 9424 7004 9470
rect 7056 9424 7070 9476
rect 6870 9420 7070 9424
rect 6990 9410 7070 9420
rect 6870 9376 7070 9380
rect 6870 9324 6884 9376
rect 6936 9324 7070 9376
rect 6870 9320 7070 9324
rect 6870 9310 6950 9320
rect 6990 9286 7070 9290
rect 6990 9280 7004 9286
rect 6870 9234 7004 9280
rect 7056 9234 7070 9286
rect 6870 9230 7070 9234
rect 6990 9220 7070 9230
rect 6870 9186 6950 9190
rect 6870 9134 6884 9186
rect 6936 9180 6950 9186
rect 6936 9134 7070 9180
rect 6870 9130 7070 9134
rect 6870 9120 6950 9130
rect 6870 9086 7070 9090
rect 6870 9040 7004 9086
rect 6990 9034 7004 9040
rect 7056 9034 7070 9086
rect 6990 9020 7070 9034
rect 6870 8996 6950 9000
rect 6870 8944 6884 8996
rect 6936 8990 6950 8996
rect 6936 8944 7070 8990
rect 6870 8940 7070 8944
rect 6870 8930 6950 8940
rect 6870 8896 7070 8900
rect 6870 8850 7004 8896
rect 6990 8844 7004 8850
rect 7056 8844 7070 8896
rect 6990 8830 7070 8844
rect 6870 8806 6950 8810
rect 6870 8754 6884 8806
rect 6936 8800 6950 8806
rect 6936 8754 7070 8800
rect 6870 8750 7070 8754
rect 6870 8740 6950 8750
rect 6990 8706 7070 8710
rect 6990 8700 7004 8706
rect 6870 8654 7004 8700
rect 7056 8654 7070 8706
rect 6870 8650 7070 8654
rect 6990 8640 7070 8650
rect 6870 8606 7070 8610
rect 6870 8554 6884 8606
rect 6936 8560 7070 8606
rect 6936 8554 6950 8560
rect 6870 8540 6950 8554
rect 6870 8506 7070 8510
rect 6870 8460 7004 8506
rect 6990 8454 7004 8460
rect 7056 8454 7070 8506
rect 6990 8440 7070 8454
rect 7100 8400 7160 9680
rect 7420 8400 7860 8420
rect 6780 8391 7860 8400
rect 6780 8340 7454 8391
rect 7420 8339 7454 8340
rect 7506 8339 7518 8391
rect 7570 8339 7582 8391
rect 7634 8339 7646 8391
rect 7698 8339 7710 8391
rect 7762 8339 7774 8391
rect 7826 8339 7860 8391
rect 7420 8310 7860 8339
rect 5720 998 6380 1040
rect 5720 562 5768 998
rect 6332 562 6380 998
rect 5720 520 6380 562
<< via1 >>
rect 5800 9429 6300 9801
rect 7004 9614 7056 9666
rect 6884 9514 6936 9566
rect 7004 9424 7056 9476
rect 6884 9324 6936 9376
rect 7004 9234 7056 9286
rect 6884 9134 6936 9186
rect 7004 9034 7056 9086
rect 6884 8944 6936 8996
rect 7004 8844 7056 8896
rect 6884 8754 6936 8806
rect 7004 8654 7056 8706
rect 6884 8554 6936 8606
rect 7004 8454 7056 8506
rect 7454 8339 7506 8391
rect 7518 8339 7570 8391
rect 7582 8339 7634 8391
rect 7646 8339 7698 8391
rect 7710 8339 7762 8391
rect 7774 8339 7826 8391
rect 5768 562 6332 998
<< metal2 >>
rect 5600 9801 6950 9830
rect 5600 9429 5800 9801
rect 6300 9566 6950 9801
rect 6300 9514 6884 9566
rect 6936 9514 6950 9566
rect 6300 9429 6950 9514
rect 5600 9400 6950 9429
rect 6650 9376 6950 9400
rect 6650 9324 6884 9376
rect 6936 9324 6950 9376
rect 6650 9186 6950 9324
rect 6650 9134 6884 9186
rect 6936 9134 6950 9186
rect 6650 8996 6950 9134
rect 6650 8944 6884 8996
rect 6936 8944 6950 8996
rect 6650 8806 6950 8944
rect 6650 8754 6884 8806
rect 6936 8754 6950 8806
rect 6650 8606 6950 8754
rect 6650 8554 6884 8606
rect 6936 8554 6950 8606
rect 6650 8430 6950 8554
rect 6990 9666 7280 9990
rect 6990 9614 7004 9666
rect 7056 9614 7280 9666
rect 6990 9476 7280 9614
rect 6990 9424 7004 9476
rect 7056 9424 7280 9476
rect 6990 9286 7280 9424
rect 6990 9234 7004 9286
rect 7056 9234 7280 9286
rect 6990 9086 7280 9234
rect 6990 9034 7004 9086
rect 7056 9034 7280 9086
rect 6990 8896 7280 9034
rect 6990 8844 7004 8896
rect 7056 8844 7280 8896
rect 6990 8706 7280 8844
rect 6990 8654 7004 8706
rect 7056 8654 7280 8706
rect 6990 8506 7280 8654
rect 6990 8454 7004 8506
rect 7056 8454 7280 8506
rect 6990 8430 7280 8454
rect 7420 8393 7860 8420
rect 7420 8391 7492 8393
rect 7548 8391 7572 8393
rect 7628 8391 7652 8393
rect 7708 8391 7732 8393
rect 7788 8391 7860 8393
rect 7420 8339 7454 8391
rect 7570 8339 7572 8391
rect 7634 8339 7646 8391
rect 7708 8339 7710 8391
rect 7826 8339 7860 8391
rect 7420 8337 7492 8339
rect 7548 8337 7572 8339
rect 7628 8337 7652 8339
rect 7708 8337 7732 8339
rect 7788 8337 7860 8339
rect 7420 8310 7860 8337
rect 5600 998 6380 1040
rect 5600 562 5768 998
rect 6332 562 6380 998
rect 5600 400 6380 562
<< via2 >>
rect 7492 8391 7548 8393
rect 7572 8391 7628 8393
rect 7652 8391 7708 8393
rect 7732 8391 7788 8393
rect 7492 8339 7506 8391
rect 7506 8339 7518 8391
rect 7518 8339 7548 8391
rect 7572 8339 7582 8391
rect 7582 8339 7628 8391
rect 7652 8339 7698 8391
rect 7698 8339 7708 8391
rect 7732 8339 7762 8391
rect 7762 8339 7774 8391
rect 7774 8339 7788 8391
rect 7492 8337 7548 8339
rect 7572 8337 7628 8339
rect 7652 8337 7708 8339
rect 7732 8337 7788 8339
rect 5782 592 6318 968
<< metal3 >>
rect 7440 8393 7840 9990
rect 7440 8337 7492 8393
rect 7548 8337 7572 8393
rect 7628 8337 7652 8393
rect 7708 8337 7732 8393
rect 7788 8337 7840 8393
rect 7440 6912 7840 8337
rect 7440 6768 7488 6912
rect 7792 6768 7840 6912
rect 7440 6740 7840 6768
rect 5720 968 6660 1040
rect 5720 592 5782 968
rect 6318 592 6660 968
rect 5720 520 6660 592
<< via3 >>
rect 7488 6768 7792 6912
<< metal4 >>
rect 7440 6912 7840 6940
rect 7440 6768 7488 6912
rect 7792 6768 7840 6912
rect 7440 6080 7840 6768
use sky130_fd_pr__cap_mim_m3_1_4RCNTW  XC2
timestamp 1663011646
transform 1 0 8750 0 1 3500
box -2150 -3100 2149 3100
use sky130_fd_pr__nfet_01v8_lvt_6BNFGK  XM41
timestamp 1663011646
transform 0 1 6970 -1 0 9063
box -733 -300 733 300
use sky130_fd_pr__res_high_po_2p85_MXEQGY  XR21
timestamp 1663011646
transform 1 0 6051 0 1 5198
box -441 -4788 441 4788
<< labels >>
rlabel metal2 s 5600 400 5760 1040 4 GND
port 1 nsew
rlabel metal2 s 5600 9400 5780 9830 4 VOP
port 2 nsew
rlabel metal2 s 6990 9680 7280 9990 4 VDD
port 3 nsew
rlabel metal3 s 7440 8410 7840 9990 4 IN
port 4 nsew
rlabel locali s 6430 8350 6730 8390 4 SUB
port 5 nsew
<< end >>
