magic
tech sky130A
magscale 1 2
timestamp 1666262531
<< error_s >>
rect -2243 -2874 -2230 -2626
rect -1995 -3088 -1982 -2874
rect -4470 -3810 7062 -3806
rect -4470 -5140 7062 -5048
<< nwell >>
rect -8726 10225 -8100 11452
<< locali >>
rect -6920 9900 -6780 10760
rect -1960 10660 4480 10940
rect -1960 10600 1560 10660
rect -2980 8990 -2820 9120
rect -3350 8950 -1990 8990
rect -7740 8580 -7620 8860
rect -3330 8480 -2030 8490
rect -3350 8450 -1960 8480
rect -9000 8140 -8880 8440
rect -14000 7490 -13900 8080
rect -10900 7490 -10800 8080
rect -14030 7480 -10800 7490
rect -860 6400 -660 6820
rect 440 6400 640 6820
rect 1720 6400 1920 6820
rect 3020 6400 3220 6820
rect 4300 6400 4400 6860
rect 4620 360 5080 400
rect 4620 200 4660 360
rect 5040 200 5080 360
rect 4620 180 5080 200
rect 4640 -40 9260 20
rect 4640 -220 9260 -160
rect 4640 -580 9260 -520
rect 4640 -960 6220 -900
rect 7680 -960 9260 -900
rect 4640 -1140 6220 -1080
rect 7740 -1140 9260 -1080
rect 4640 -1500 6220 -1440
rect 7580 -1480 9260 -1420
rect 4640 -1880 9260 -1820
rect 4640 -2060 9260 -2000
rect -1860 -2560 -1560 -2400
rect -1440 -2440 4360 -2400
rect 4640 -2420 9260 -2360
rect -1440 -2460 4460 -2440
rect -1440 -2520 4520 -2460
rect -1440 -2560 4400 -2520
rect -1860 -2580 4400 -2560
rect 4300 -2780 4400 -2580
rect 8480 -2780 9420 -2740
rect 7700 -3420 9500 -3260
rect -14180 -3820 -13640 -3520
rect 7700 -3960 9500 -3840
rect -14200 -10160 -13640 -9020
rect 8100 -10296 9500 -10200
<< viali >>
rect -10880 10080 -10820 11240
rect -8800 10200 -8680 10580
rect -2980 9120 -2820 9280
rect 4660 200 5040 360
rect -1560 -2560 -1440 -2400
rect 9620 -2960 9920 -2840
rect 33500 -2960 33800 -2840
rect 61800 -2960 62100 -2840
<< metal1 >>
rect -10910 10060 -10900 11260
rect -10800 10060 -10790 11260
rect -7750 11040 -7740 11120
rect -7680 11040 -7670 11120
rect 1190 11100 1200 11200
rect 1300 11100 1310 11200
rect -11458 9858 -10653 9906
rect -10600 8810 -10540 11000
rect -8806 10580 -8674 10592
rect -8810 10200 -8800 10580
rect -8680 10200 -8670 10580
rect -8230 10500 -8220 10580
rect -8140 10500 -7760 10580
rect -8806 10188 -8674 10200
rect -7780 9760 -7640 9920
rect -2992 9280 -2808 9286
rect -2992 9120 -2980 9280
rect -2820 9120 -2808 9280
rect -8630 9040 -8620 9120
rect -8560 9040 -8550 9120
rect -2992 9114 -2808 9120
rect -8850 8810 -8840 8820
rect -13422 8764 -8840 8810
rect -10600 8760 -10540 8764
rect -8850 8760 -8840 8764
rect -8780 8760 -8770 8820
rect -7950 8760 -7940 8820
rect -7880 8760 -7870 8820
rect -8700 8200 -4700 8400
rect -10090 7800 -10080 7860
rect -10020 7800 -9100 7860
rect -9200 5800 -9100 7800
rect -8710 6000 -8700 6100
rect -8600 6000 -8590 6100
rect -13300 5700 -9100 5800
rect -13300 5020 -13200 5700
rect -9200 -100 -9100 5700
rect -4900 4000 -4700 8200
rect -4900 3800 -700 4000
rect 4648 360 5052 366
rect 4648 200 4660 360
rect 5040 200 5052 360
rect 4648 194 5052 200
rect -13300 -200 -9100 -100
rect -13300 -900 -13200 -200
rect -9200 -3200 -9100 -200
rect 6180 -1220 6980 -1160
rect -1566 -2400 -1434 -2388
rect -1570 -2560 -1560 -2400
rect -1440 -2560 -1430 -2400
rect -1566 -2572 -1434 -2560
rect -1770 -3060 -1760 -2940
rect -1660 -3060 -1650 -2940
rect 6180 -3480 6260 -1220
rect 9608 -2840 9932 -2834
rect 9608 -2960 9620 -2840
rect 9920 -2960 9932 -2840
rect 8110 -3060 8120 -2960
rect 8200 -3060 8210 -2960
rect 9608 -2966 9932 -2960
rect 33488 -2840 33812 -2834
rect 33488 -2960 33500 -2840
rect 33800 -2960 33812 -2840
rect 33488 -2966 33812 -2960
rect 61788 -2840 62112 -2834
rect 61788 -2960 61800 -2840
rect 62100 -2960 62112 -2840
rect 61788 -2966 62112 -2960
rect 6080 -3540 6360 -3480
rect -14180 -3560 -13640 -3540
rect -14180 -3780 -14140 -3560
rect -13660 -3780 -13640 -3560
rect 6140 -3660 6360 -3540
rect 6080 -3700 6360 -3660
rect 6600 -3540 7600 -3500
rect 6600 -3660 6640 -3540
rect 6720 -3660 7600 -3540
rect 6600 -3700 7600 -3660
rect -14180 -3800 -13640 -3780
rect -11660 -3820 7040 -3800
rect -11660 -3860 6940 -3820
rect -11660 -3960 -11500 -3860
rect -11400 -3960 6940 -3860
rect 7020 -3960 7040 -3820
rect -11660 -4000 7040 -3960
rect 6800 -4500 7040 -4000
rect 6800 -4700 7800 -4500
rect -14200 -9200 -13640 -9020
rect -14200 -10000 -14100 -9200
rect -13700 -10000 -13640 -9200
rect -14200 -10160 -13640 -10000
rect 9590 -10360 9600 -10240
rect 9900 -10360 9910 -10240
rect 35690 -10360 35700 -10240
rect 35996 -10360 36006 -10240
rect 61790 -10360 61800 -10240
rect 62100 -10360 62110 -10240
<< via1 >>
rect -10900 11240 -10800 11260
rect -10900 10080 -10880 11240
rect -10880 10080 -10820 11240
rect -10820 10080 -10800 11240
rect -10900 10060 -10800 10080
rect -7740 11040 -7680 11120
rect 1200 11100 1300 11200
rect -8800 10200 -8680 10580
rect -8220 10500 -8140 10580
rect -2980 9120 -2820 9280
rect -8620 9040 -8560 9120
rect -8840 8760 -8780 8820
rect -7940 8760 -7880 8820
rect -10080 7800 -10020 7860
rect -8700 6000 -8600 6100
rect 4660 200 5040 360
rect -1560 -2560 -1440 -2400
rect -1760 -3060 -1660 -2940
rect 9620 -2960 9920 -2840
rect 8120 -3060 8200 -2960
rect 33500 -2960 33800 -2840
rect 61800 -2960 62100 -2840
rect -14140 -3780 -13660 -3560
rect 6080 -3660 6140 -3540
rect 6640 -3660 6720 -3540
rect -11500 -3960 -11400 -3860
rect 6940 -3960 7020 -3820
rect -14100 -10000 -13700 -9200
rect 9600 -10360 9900 -10240
rect 35700 -10360 35996 -10240
rect 61800 -10360 62100 -10240
<< metal2 >>
rect -10900 11260 -10800 11270
rect -10800 11186 -10642 11246
rect -7900 11140 -7700 12500
rect 1160 11200 1380 11220
rect -8940 11120 -7680 11140
rect -8940 11040 -7740 11120
rect -8940 11020 -7680 11040
rect 1160 11100 1200 11200
rect 1300 11100 1380 11200
rect -10800 10826 -10648 10886
rect -8480 10860 -8400 10870
rect -8800 10580 -8680 10590
rect -10800 10446 -10656 10506
rect -8800 10190 -8680 10200
rect -10800 10086 -10650 10146
rect -10900 9680 -10800 10060
rect -9100 9780 -9000 10000
rect -9100 9720 -9080 9780
rect -9020 9720 -9000 9780
rect -9100 9700 -9000 9720
rect -10900 9620 -10620 9680
rect -10900 9320 -10800 9620
rect -8660 9520 -8600 9530
rect -9440 9460 -8660 9520
rect -8660 9450 -8600 9460
rect -10900 9260 -10620 9320
rect -10900 9240 -10800 9260
rect -14160 8460 -13540 8520
rect -14160 5760 -14100 8460
rect -11260 7680 -11180 8700
rect -10080 7860 -10020 9160
rect -8620 9120 -8560 9130
rect -8480 9120 -8400 10780
rect -8220 10580 -8140 10590
rect -8220 10490 -8140 10500
rect -8560 9040 -8400 9120
rect -2980 9280 -2820 9290
rect -2980 9110 -2820 9120
rect -8620 9030 -8560 9040
rect -8860 8840 -8760 8850
rect -8860 8730 -8760 8740
rect -8216 8840 -8114 8940
rect -8216 8820 -7880 8840
rect -8216 8760 -8200 8820
rect -8140 8760 -7940 8820
rect 1160 8800 1380 11100
rect -8216 8740 -7880 8760
rect -10080 7790 -10020 7800
rect -11260 7620 -9480 7680
rect -9540 6100 -9480 7620
rect -8216 6980 -8114 8740
rect 1200 8700 1300 8800
rect -8700 6100 -8600 6110
rect -9540 6000 -8700 6100
rect -11600 5760 -11540 5770
rect -14160 5700 -11600 5760
rect -11600 5690 -11540 5700
rect -11460 5760 -11400 5770
rect -9540 5760 -9480 6000
rect -8700 5990 -8600 6000
rect -11400 5700 -9480 5760
rect -11460 5690 -11400 5700
rect -11460 5120 -11400 5130
rect -11460 4280 -11400 5060
rect 6400 4400 28300 4600
rect -11520 4240 -11400 4280
rect -11620 4100 -11500 4126
rect -11620 4040 -11600 4100
rect -11540 4040 -11500 4100
rect -11620 4000 -11500 4040
rect -11280 3180 -11220 3190
rect -11280 2500 -11220 3120
rect -11280 2300 1300 2500
rect 1060 1820 1300 2300
rect 4660 360 5040 370
rect 6420 320 6600 4400
rect 28000 4300 28300 4400
rect 27200 4100 29100 4300
rect 29400 4260 31300 4300
rect 29400 4140 30240 4260
rect 30460 4140 31300 4260
rect 29400 4100 31300 4140
rect 31600 4260 33500 4300
rect 31600 4140 32440 4260
rect 32660 4140 33500 4260
rect 31600 4100 33500 4140
rect 33800 4260 35700 4300
rect 33800 4140 34640 4260
rect 34860 4140 35700 4260
rect 33800 4100 35700 4140
rect 36000 4260 37900 4300
rect 36000 4140 36840 4260
rect 37060 4140 37900 4260
rect 36000 4100 37900 4140
rect 38200 4260 40100 4300
rect 38200 4140 39040 4260
rect 39260 4140 40100 4260
rect 38200 4100 40100 4140
rect 40400 4260 42300 4300
rect 40400 4140 41240 4260
rect 41460 4140 42300 4260
rect 40400 4100 42300 4140
rect 42600 4260 44500 4300
rect 42600 4140 43440 4260
rect 43660 4140 44500 4260
rect 42600 4100 44500 4140
rect 6420 240 6480 320
rect 6540 240 6600 320
rect 6480 230 6540 240
rect 4660 190 5040 200
rect 6460 -840 6660 -820
rect 6540 -940 6660 -840
rect 6460 -960 6660 -940
rect 6900 -1460 7180 -1380
rect 6900 -1540 6920 -1460
rect 7040 -1540 7180 -1460
rect 6900 -1560 7180 -1540
rect -11540 -1620 -11420 -1600
rect -11540 -1680 -11520 -1620
rect -11440 -1680 -11420 -1620
rect -11540 -1700 -11420 -1680
rect -11880 -1800 -11780 -1790
rect -11880 -1890 -11780 -1880
rect -1560 -2400 -1440 -2390
rect -1560 -2570 -1440 -2560
rect 28000 -2800 28300 -2600
rect 9620 -2840 9920 -2830
rect -1800 -2940 6720 -2900
rect -5600 -3500 -5400 -3000
rect -1800 -3060 -1760 -2940
rect -1660 -3060 6720 -2940
rect -1800 -3100 6720 -3060
rect 6920 -2960 8240 -2940
rect 6920 -3060 6940 -2960
rect 7020 -3060 8120 -2960
rect 8200 -3060 8240 -2960
rect 28000 -2880 28040 -2800
rect 28260 -2880 28300 -2800
rect 28000 -2900 28300 -2880
rect 30200 -2800 30500 -2600
rect 30200 -2880 30240 -2800
rect 30460 -2880 30500 -2800
rect 30200 -2900 30500 -2880
rect 32400 -2800 32700 -2600
rect 32400 -2880 32440 -2800
rect 32660 -2880 32700 -2800
rect 34600 -2800 34900 -2600
rect 32400 -2900 32700 -2880
rect 33500 -2840 33800 -2830
rect 9620 -2970 9920 -2960
rect 34600 -2880 34640 -2800
rect 34860 -2880 34900 -2800
rect 34600 -2900 34900 -2880
rect 36800 -2800 37100 -2600
rect 36800 -2880 36840 -2800
rect 37060 -2880 37100 -2800
rect 36800 -2900 37100 -2880
rect 39000 -2800 39300 -2600
rect 39000 -2880 39040 -2800
rect 39260 -2880 39300 -2800
rect 39000 -2900 39300 -2880
rect 41200 -2800 41500 -2600
rect 41200 -2880 41240 -2800
rect 41460 -2880 41500 -2800
rect 41200 -2900 41500 -2880
rect 43400 -2800 43700 -2600
rect 43400 -2880 43440 -2800
rect 43660 -2880 43700 -2800
rect 43400 -2900 43700 -2880
rect 61800 -2840 62100 -2830
rect 33500 -2970 33800 -2960
rect 61800 -2970 62100 -2960
rect 6920 -3080 8240 -3060
rect 5980 -3500 6360 -3480
rect -5600 -3540 6360 -3500
rect -14140 -3560 -13660 -3550
rect -5600 -3660 6080 -3540
rect 6140 -3660 6360 -3540
rect -5600 -3700 6360 -3660
rect 6600 -3540 6720 -3100
rect 6600 -3660 6640 -3540
rect 6600 -3680 6720 -3660
rect -14140 -3790 -13660 -3780
rect 6940 -3800 7020 -3790
rect -11500 -3860 -11400 -3850
rect -11500 -3970 -11400 -3960
rect 6940 -3990 7020 -3980
rect -14100 -9200 -13700 -9190
rect -14100 -10010 -13700 -10000
rect 9600 -10240 9900 -10230
rect 9600 -10370 9900 -10360
rect 35700 -10240 35996 -10230
rect 35700 -10370 35996 -10360
rect 61800 -10240 62100 -10230
rect 61800 -10370 62100 -10360
<< via2 >>
rect -10900 10060 -10800 11260
rect -8480 10780 -8400 10860
rect -8800 10200 -8680 10580
rect -9080 9720 -9020 9780
rect -8660 9460 -8600 9520
rect -8220 10500 -8140 10580
rect -2980 9120 -2820 9280
rect -8860 8820 -8760 8840
rect -8860 8760 -8840 8820
rect -8840 8760 -8780 8820
rect -8780 8760 -8760 8820
rect -8860 8740 -8760 8760
rect -8200 8760 -8140 8820
rect -11600 5700 -11540 5760
rect -11460 5700 -11400 5760
rect -11460 5060 -11400 5120
rect -11600 4040 -11540 4100
rect -11280 3120 -11220 3180
rect 4660 200 5040 360
rect 30240 4140 30460 4260
rect 32440 4140 32660 4260
rect 34640 4140 34860 4260
rect 36840 4140 37060 4260
rect 39040 4140 39260 4260
rect 41240 4140 41460 4260
rect 43440 4140 43660 4260
rect 6480 240 6540 320
rect 6460 -940 6540 -840
rect 6920 -1540 7040 -1460
rect -11520 -1680 -11440 -1620
rect -11880 -1880 -11780 -1800
rect -1560 -2560 -1440 -2400
rect 6940 -3060 7020 -2960
rect 9620 -2960 9920 -2840
rect 28040 -2880 28260 -2800
rect 30240 -2880 30460 -2800
rect 32440 -2880 32660 -2800
rect 33500 -2960 33800 -2840
rect 34640 -2880 34860 -2800
rect 36840 -2880 37060 -2800
rect 39040 -2880 39260 -2800
rect 41240 -2880 41460 -2800
rect 43440 -2880 43660 -2800
rect 61800 -2960 62100 -2840
rect -14140 -3780 -13660 -3560
rect 6940 -3820 7020 -3800
rect -11500 -3960 -11400 -3860
rect 6940 -3960 7020 -3820
rect 6940 -3980 7020 -3960
rect -14100 -10000 -13700 -9200
rect 9600 -10360 9900 -10240
rect 35700 -10360 35996 -10240
rect 61800 -10360 62100 -10240
<< metal3 >>
rect -10910 11260 -10790 11265
rect -10910 10060 -10900 11260
rect -10800 10060 -10790 11260
rect -8500 10860 -8380 12540
rect -8500 10780 -8480 10860
rect -8400 10780 -8380 10860
rect -8500 10760 -8380 10780
rect -8810 10580 -8670 10585
rect -8810 10200 -8800 10580
rect -8680 10200 -8670 10580
rect -8230 10580 -8130 10585
rect -8230 10500 -8220 10580
rect -8140 10500 -8130 10580
rect -8230 10495 -8130 10500
rect -8810 10195 -8670 10200
rect -10910 10055 -10790 10060
rect -9100 9780 -9000 9800
rect -14190 9726 -14180 9760
rect -14200 9666 -14180 9726
rect -14190 9620 -14180 9666
rect -14060 9726 -14050 9760
rect -10910 9726 -10900 9740
rect -14060 9666 -13460 9726
rect -11340 9666 -10900 9726
rect -14060 9620 -14050 9666
rect -10910 9640 -10900 9666
rect -10800 9640 -10790 9740
rect -9100 9720 -9080 9780
rect -9020 9720 -9000 9780
rect -11610 5760 -11530 5790
rect -11610 5700 -11600 5760
rect -11540 5700 -11530 5760
rect -11610 4100 -11530 5700
rect -11470 5760 -11390 5770
rect -11470 5700 -11460 5760
rect -11400 5700 -11390 5760
rect -11470 5120 -11390 5700
rect -11470 5060 -11460 5120
rect -11400 5060 -11390 5120
rect -11470 5050 -11390 5060
rect -11610 4040 -11600 4100
rect -11540 4040 -11530 4100
rect -11610 3200 -11530 4040
rect -11610 3180 -11200 3200
rect -11610 3120 -11280 3180
rect -11220 3120 -11200 3180
rect -11290 3115 -11210 3120
rect -9100 2200 -9000 9720
rect -8220 9540 -8140 10495
rect -8680 9520 -8140 9540
rect -8680 9460 -8660 9520
rect -8600 9460 -8140 9520
rect -8680 9440 -8140 9460
rect -2990 9280 -2810 9285
rect -2990 9120 -2980 9280
rect -2820 9120 -2810 9280
rect -2990 9115 -2810 9120
rect -8870 8840 -8750 8845
rect -8870 8740 -8860 8840
rect -8760 8820 -8120 8840
rect -8760 8760 -8200 8820
rect -8140 8760 -8120 8820
rect -8760 8740 -8120 8760
rect -8870 8735 -8750 8740
rect 30200 4260 30500 12600
rect 30200 4140 30240 4260
rect 30460 4140 30500 4260
rect 30200 4100 30500 4140
rect 32400 4260 32700 12600
rect 32400 4140 32440 4260
rect 32660 4140 32700 4260
rect 32400 4100 32700 4140
rect 34600 4260 34900 12600
rect 34600 4140 34640 4260
rect 34860 4140 34900 4260
rect 34600 4100 34900 4140
rect 36800 4260 37100 12600
rect 36800 4140 36840 4260
rect 37060 4140 37100 4260
rect 36800 4100 37100 4140
rect 39000 4260 39300 12600
rect 39000 4140 39040 4260
rect 39260 4140 39300 4260
rect 39000 4100 39300 4140
rect 41200 4260 41500 12600
rect 41200 4140 41240 4260
rect 41460 4140 41500 4260
rect 41200 4100 41500 4140
rect 43400 4260 43700 12600
rect 43400 4140 43440 4260
rect 43660 4140 43700 4260
rect 43400 4100 43700 4140
rect -7040 3240 -6880 4060
rect -7040 3040 -7020 3240
rect -6900 3040 -6880 3240
rect -7040 2200 -6880 3040
rect -11900 2100 -9000 2200
rect -11900 -1795 -11800 2100
rect 4650 360 5050 365
rect 4650 200 4660 360
rect 5040 200 5050 360
rect 4650 195 5050 200
rect 6460 320 6560 340
rect 6460 240 6480 320
rect 6540 240 6560 320
rect 6460 -835 6560 240
rect 6450 -840 6560 -835
rect 6450 -940 6460 -840
rect 6540 -940 6560 -840
rect 6450 -945 6550 -940
rect 6910 -1460 7050 -1455
rect 6910 -1540 6920 -1460
rect 7040 -1540 7050 -1460
rect 6910 -1545 7050 -1540
rect -11480 -1615 -11420 -1600
rect -11530 -1620 -11420 -1615
rect -11530 -1680 -11520 -1620
rect -11440 -1680 -11420 -1620
rect -11530 -1685 -11420 -1680
rect -11900 -1800 -11770 -1795
rect -11900 -1880 -11880 -1800
rect -11780 -1880 -11770 -1800
rect -11900 -1885 -11770 -1880
rect -11900 -1900 -11800 -1885
rect -14150 -3560 -13650 -3555
rect -14150 -3780 -14140 -3560
rect -13660 -3780 -13650 -3560
rect -14150 -3785 -13650 -3780
rect -11480 -3855 -11420 -1685
rect -1570 -2400 -1430 -2395
rect -1570 -2560 -1560 -2400
rect -1440 -2560 -1430 -2400
rect -1570 -2565 -1430 -2560
rect 6920 -2960 7040 -1545
rect 28030 -2800 28270 -2795
rect 6920 -3060 6940 -2960
rect 7020 -3060 7040 -2960
rect 9610 -2840 9930 -2835
rect 9610 -2960 9620 -2840
rect 9920 -2960 9930 -2840
rect 28030 -2880 28040 -2800
rect 28260 -2880 28270 -2800
rect 28030 -2885 28270 -2880
rect 30230 -2800 30470 -2795
rect 30230 -2880 30240 -2800
rect 30460 -2880 30470 -2800
rect 30230 -2885 30470 -2880
rect 32430 -2800 32670 -2795
rect 32430 -2880 32440 -2800
rect 32660 -2880 32670 -2800
rect 34630 -2800 34870 -2795
rect 32430 -2885 32670 -2880
rect 33490 -2840 33810 -2835
rect 9610 -2965 9930 -2960
rect 33490 -2960 33500 -2840
rect 33800 -2960 33810 -2840
rect 34630 -2880 34640 -2800
rect 34860 -2880 34870 -2800
rect 34630 -2885 34870 -2880
rect 36830 -2800 37070 -2795
rect 36830 -2880 36840 -2800
rect 37060 -2880 37070 -2800
rect 36830 -2885 37070 -2880
rect 39030 -2800 39270 -2795
rect 39030 -2880 39040 -2800
rect 39260 -2880 39270 -2800
rect 39030 -2885 39270 -2880
rect 41230 -2800 41470 -2795
rect 41230 -2880 41240 -2800
rect 41460 -2880 41470 -2800
rect 41230 -2885 41470 -2880
rect 43430 -2800 43670 -2795
rect 43430 -2880 43440 -2800
rect 43660 -2880 43670 -2800
rect 43430 -2885 43670 -2880
rect 61790 -2840 62110 -2835
rect 33490 -2965 33810 -2960
rect 61790 -2960 61800 -2840
rect 62100 -2960 62110 -2840
rect 61790 -2965 62110 -2960
rect 6920 -3800 7040 -3060
rect -11510 -3860 -11390 -3855
rect -11510 -3960 -11500 -3860
rect -11400 -3960 -11390 -3860
rect -11510 -3965 -11390 -3960
rect 6920 -3980 6940 -3800
rect 7020 -3980 7040 -3800
rect 6920 -4000 7040 -3980
rect -14110 -9200 -13690 -9195
rect -14110 -10000 -14100 -9200
rect -13700 -10000 -13690 -9200
rect -14110 -10005 -13690 -10000
rect 9590 -10240 9910 -10235
rect 9590 -10360 9600 -10240
rect 9900 -10360 9910 -10240
rect 9590 -10365 9910 -10360
rect 35690 -10240 36006 -10235
rect 35690 -10360 35700 -10240
rect 35996 -10360 36006 -10240
rect 35690 -10365 36006 -10360
rect 61790 -10240 62110 -10235
rect 61790 -10360 61800 -10240
rect 62100 -10360 62110 -10240
rect 61790 -10365 62110 -10360
<< via3 >>
rect -10900 10060 -10800 11260
rect -8800 10200 -8680 10580
rect -14180 9620 -14060 9760
rect -10900 9640 -10800 9740
rect -2980 9120 -2820 9280
rect -7020 3040 -6900 3240
rect 4660 200 5040 360
rect -14140 -3780 -13660 -3560
rect -1560 -2560 -1440 -2400
rect 9620 -2960 9920 -2840
rect 28040 -2880 28260 -2800
rect 30240 -2880 30460 -2800
rect 32440 -2880 32660 -2800
rect 33500 -2960 33800 -2840
rect 34640 -2880 34860 -2800
rect 36840 -2880 37060 -2800
rect 39040 -2880 39260 -2800
rect 41240 -2880 41460 -2800
rect 43440 -2880 43660 -2800
rect 61800 -2960 62100 -2840
rect -14100 -10000 -13700 -9200
rect 9600 -10360 9900 -10240
rect 35700 -10360 35996 -10240
rect 61800 -10360 62100 -10240
<< metal4 >>
rect -14220 11800 62300 12000
rect -14220 9760 -14020 11800
rect -14220 9620 -14180 9760
rect -14060 9620 -14020 9760
rect -14220 7400 -14020 9620
rect -10920 11260 -10780 11800
rect -10920 10060 -10900 11260
rect -10800 10060 -10780 11260
rect -8800 10581 -8600 11800
rect -8801 10580 -8600 10581
rect -8801 10200 -8800 10580
rect -8680 10200 -8600 10580
rect -8801 10199 -8600 10200
rect -10920 9740 -10780 10060
rect -10920 9640 -10900 9740
rect -10800 9640 -10780 9740
rect -10920 7580 -10780 9640
rect -8800 7500 -8600 10199
rect -3500 9280 -2800 9300
rect -3500 9120 -2980 9280
rect -2820 9120 -2800 9280
rect -3500 9100 -2800 9120
rect -7021 3240 -6899 3241
rect 4600 3240 4800 11800
rect -7021 3040 -7020 3240
rect -6900 3040 4800 3240
rect -7021 3039 -6899 3040
rect -2140 2540 -1400 2740
rect -1600 -2400 -1400 2540
rect 4600 400 4800 3040
rect 4600 360 5100 400
rect 4600 200 4660 360
rect 5040 200 5100 360
rect 4600 180 5100 200
rect -1600 -2560 -1560 -2400
rect -1440 -2560 -1400 -2400
rect -1600 -3180 -1400 -2560
rect 28039 -2800 28261 -2799
rect 30239 -2800 30461 -2799
rect 32439 -2800 32661 -2799
rect 34639 -2800 34861 -2799
rect 36839 -2800 37061 -2799
rect 39039 -2800 39261 -2799
rect 41239 -2800 41461 -2799
rect 43439 -2800 43661 -2799
rect 9300 -2840 28040 -2800
rect 9300 -2960 9620 -2840
rect 9920 -2880 28040 -2840
rect 28260 -2880 30240 -2800
rect 30460 -2880 32440 -2800
rect 32660 -2840 34640 -2800
rect 32660 -2880 33500 -2840
rect 9920 -2960 33500 -2880
rect 33800 -2880 34640 -2840
rect 34860 -2880 36840 -2800
rect 37060 -2880 39040 -2800
rect 39260 -2880 41240 -2800
rect 41460 -2880 43440 -2800
rect 43660 -2840 62400 -2800
rect 43660 -2880 61800 -2840
rect 33800 -2960 61800 -2880
rect 62100 -2960 62400 -2840
rect 9300 -3000 62400 -2960
rect -14220 -3559 -14020 -3240
rect -2580 -3380 -1380 -3180
rect -1600 -3400 -1400 -3380
rect -14220 -3560 -13659 -3559
rect -14220 -3780 -14140 -3560
rect -13660 -3780 -13659 -3560
rect -14220 -3781 -13659 -3780
rect -14220 -9199 -14020 -3781
rect -14220 -9200 -13699 -9199
rect -14220 -10000 -14100 -9200
rect -13700 -10000 -13699 -9200
rect -14220 -10001 -13699 -10000
rect -14220 -10200 -14020 -10001
rect 9300 -10200 9600 -3000
rect 62200 -10200 62400 -3000
rect -14220 -10240 62400 -10200
rect -14220 -10360 9600 -10240
rect 9900 -10360 35700 -10240
rect 35996 -10360 61800 -10240
rect 62100 -10360 62400 -10240
rect -14220 -10400 62400 -10360
use XM_Rref  XM_Rref_0
timestamp 1665771957
transform 0 1 -13057 -1 0 -5305
box -1417 -1173 5029 21223
use XM_bjt  XM_bjt_0
timestamp 1666262531
transform 1 0 -1950 0 1 -2620
box 0 0 6492 9068
use XM_bjt_out  XM_bjt_out_0
timestamp 1666262531
transform 1 0 -2070 0 1 6780
box 0 0 6492 3916
use XM_current_gate_with_dummy  XM_current_gate_with_dummy_0
timestamp 1662842659
transform 1 0 4644 0 1 -1712
box 0 -924 4660 1954
use XM_feedbackmir2  XM_feedbackmir2_0
timestamp 1662719914
transform 1 0 -10768 0 1 9846
box -140 -160 2080 1600
use XM_feedbackmir  XM_feedbackmir_0
timestamp 1662675866
transform 1 0 -13500 0 1 8386
box -700 -500 2900 3100
use XM_otabias_nmos  XM_otabias_nmos_0
timestamp 1662916051
transform 1 0 -7877 0 1 9671
box -53 -53 1139 1305
use XM_otabias_pmos  XM_otabias_pmos_0
timestamp 1662818872
transform 1 0 -10817 0 1 8939
box -53 -53 1571 879
use XM_output_mirr_combined_with_dummy  XM_output_mirr_combined_with_dummy_0
timestamp 1662903677
transform 1 0 26905 0 1 -3003
box -17600 -7400 35500 15000
use XM_pdn  XM_pdn_0
timestamp 1662820526
transform 1 0 -8785 0 1 9133
box -53 -718 5502 1206
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_0
timestamp 1662836520
transform 1 0 -8840 0 1 1874
box -5380 594 6776 6403
use opamp_realcomp3_usefinger  opamp_realcomp3_usefinger_1
timestamp 1662836520
transform 1 0 -8840 0 1 -4044
box -5380 594 6776 6403
use sky130_fd_pr__res_high_po_1p41_6ZUZ5C  sky130_fd_pr__res_high_po_1p41_6ZUZ5C_0
timestamp 1662820359
transform 1 0 -8623 0 1 7103
box -307 -1408 307 1408
use sky130_fd_pr__res_high_po_1p41_GWJZ59  sky130_fd_pr__res_high_po_1p41_GWJZ59_0
timestamp 1663020457
transform 0 1 -3232 -1 0 -3669
box -307 -10998 307 10998
use sky130_fd_pr__res_high_po_1p41_HX7ZEK  sky130_fd_pr__res_high_po_1p41_HX7ZEK_0
timestamp 1662827686
transform 0 1 3187 -1 0 -3015
box -307 -5348 307 5348
use sky130_fd_pr__res_high_po_1p41_S8KB58  sky130_fd_pr__res_high_po_1p41_S8KB58_0
timestamp 1662758895
transform 0 1 -3253 -1 0 11177
box -307 -4837 307 4837
<< labels >>
rlabel metal2 -9540 5700 -9480 7680 0 vb
rlabel metal3 -8760 8740 -8200 8840 0 vgate
rlabel metal2 1160 8800 1380 11100 0 vbe3
rlabel metal1 -9200 -2991 -9100 5271 0 Vota_bias1
rlabel space -11280 2300 1400 2500 0 va
rlabel metal3 6920 -3800 7040 -1540 0 vd4
rlabel metal2 6420 320 6600 4600 0 voutb2
rlabel space -3765 8753 -3645 10339 0 porst_buff
rlabel space 27267 -1013 29033 -859 0 voutb1
rlabel metal1 -8700 8200 -4700 8400 0 vbneg
rlabel metal3 30200 4260 30500 12600 0 Iout0
port 1 nsew
rlabel metal4 -14220 9760 -14020 12000 0 VDD
port 2 nsew
rlabel metal4 -14220 -9200 -14020 -3780 0 VSS
port 3 nsew
rlabel metal3 32400 4260 32700 12600 0 Iout1
port 4 nsew
rlabel metal3 34600 4260 34900 12600 0 Iout2
port 5 nsew
rlabel metal3 -8500 10860 -8380 12540 0 porst
port 6 nsew
rlabel metal2 -7900 11120 -7700 12500 0 vbg
port 7 nsew
rlabel metal3 36800 4260 37100 12600 0 Iout3
port 8 nsew
rlabel metal3 39000 4260 39300 12600 0 Iout4
port 9 nsew
rlabel metal3 41200 4260 41500 12600 0 Iout5
port 10 nsew
rlabel metal3 43400 4260 43700 12600 0 Iout6
port 11 nsew
<< end >>
