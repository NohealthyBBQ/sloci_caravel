magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -615 -1481 615 1481
<< nmoslvt >>
rect -429 943 -29 1343
rect 29 943 429 1343
rect -429 387 -29 787
rect 29 387 429 787
rect -429 -169 -29 231
rect 29 -169 429 231
rect -429 -725 -29 -325
rect 29 -725 429 -325
rect -429 -1281 -29 -881
rect 29 -1281 429 -881
<< ndiff >>
rect -487 1330 -429 1343
rect -487 1296 -475 1330
rect -441 1296 -429 1330
rect -487 1262 -429 1296
rect -487 1228 -475 1262
rect -441 1228 -429 1262
rect -487 1194 -429 1228
rect -487 1160 -475 1194
rect -441 1160 -429 1194
rect -487 1126 -429 1160
rect -487 1092 -475 1126
rect -441 1092 -429 1126
rect -487 1058 -429 1092
rect -487 1024 -475 1058
rect -441 1024 -429 1058
rect -487 990 -429 1024
rect -487 956 -475 990
rect -441 956 -429 990
rect -487 943 -429 956
rect -29 1330 29 1343
rect -29 1296 -17 1330
rect 17 1296 29 1330
rect -29 1262 29 1296
rect -29 1228 -17 1262
rect 17 1228 29 1262
rect -29 1194 29 1228
rect -29 1160 -17 1194
rect 17 1160 29 1194
rect -29 1126 29 1160
rect -29 1092 -17 1126
rect 17 1092 29 1126
rect -29 1058 29 1092
rect -29 1024 -17 1058
rect 17 1024 29 1058
rect -29 990 29 1024
rect -29 956 -17 990
rect 17 956 29 990
rect -29 943 29 956
rect 429 1330 487 1343
rect 429 1296 441 1330
rect 475 1296 487 1330
rect 429 1262 487 1296
rect 429 1228 441 1262
rect 475 1228 487 1262
rect 429 1194 487 1228
rect 429 1160 441 1194
rect 475 1160 487 1194
rect 429 1126 487 1160
rect 429 1092 441 1126
rect 475 1092 487 1126
rect 429 1058 487 1092
rect 429 1024 441 1058
rect 475 1024 487 1058
rect 429 990 487 1024
rect 429 956 441 990
rect 475 956 487 990
rect 429 943 487 956
rect -487 774 -429 787
rect -487 740 -475 774
rect -441 740 -429 774
rect -487 706 -429 740
rect -487 672 -475 706
rect -441 672 -429 706
rect -487 638 -429 672
rect -487 604 -475 638
rect -441 604 -429 638
rect -487 570 -429 604
rect -487 536 -475 570
rect -441 536 -429 570
rect -487 502 -429 536
rect -487 468 -475 502
rect -441 468 -429 502
rect -487 434 -429 468
rect -487 400 -475 434
rect -441 400 -429 434
rect -487 387 -429 400
rect -29 774 29 787
rect -29 740 -17 774
rect 17 740 29 774
rect -29 706 29 740
rect -29 672 -17 706
rect 17 672 29 706
rect -29 638 29 672
rect -29 604 -17 638
rect 17 604 29 638
rect -29 570 29 604
rect -29 536 -17 570
rect 17 536 29 570
rect -29 502 29 536
rect -29 468 -17 502
rect 17 468 29 502
rect -29 434 29 468
rect -29 400 -17 434
rect 17 400 29 434
rect -29 387 29 400
rect 429 774 487 787
rect 429 740 441 774
rect 475 740 487 774
rect 429 706 487 740
rect 429 672 441 706
rect 475 672 487 706
rect 429 638 487 672
rect 429 604 441 638
rect 475 604 487 638
rect 429 570 487 604
rect 429 536 441 570
rect 475 536 487 570
rect 429 502 487 536
rect 429 468 441 502
rect 475 468 487 502
rect 429 434 487 468
rect 429 400 441 434
rect 475 400 487 434
rect 429 387 487 400
rect -487 218 -429 231
rect -487 184 -475 218
rect -441 184 -429 218
rect -487 150 -429 184
rect -487 116 -475 150
rect -441 116 -429 150
rect -487 82 -429 116
rect -487 48 -475 82
rect -441 48 -429 82
rect -487 14 -429 48
rect -487 -20 -475 14
rect -441 -20 -429 14
rect -487 -54 -429 -20
rect -487 -88 -475 -54
rect -441 -88 -429 -54
rect -487 -122 -429 -88
rect -487 -156 -475 -122
rect -441 -156 -429 -122
rect -487 -169 -429 -156
rect -29 218 29 231
rect -29 184 -17 218
rect 17 184 29 218
rect -29 150 29 184
rect -29 116 -17 150
rect 17 116 29 150
rect -29 82 29 116
rect -29 48 -17 82
rect 17 48 29 82
rect -29 14 29 48
rect -29 -20 -17 14
rect 17 -20 29 14
rect -29 -54 29 -20
rect -29 -88 -17 -54
rect 17 -88 29 -54
rect -29 -122 29 -88
rect -29 -156 -17 -122
rect 17 -156 29 -122
rect -29 -169 29 -156
rect 429 218 487 231
rect 429 184 441 218
rect 475 184 487 218
rect 429 150 487 184
rect 429 116 441 150
rect 475 116 487 150
rect 429 82 487 116
rect 429 48 441 82
rect 475 48 487 82
rect 429 14 487 48
rect 429 -20 441 14
rect 475 -20 487 14
rect 429 -54 487 -20
rect 429 -88 441 -54
rect 475 -88 487 -54
rect 429 -122 487 -88
rect 429 -156 441 -122
rect 475 -156 487 -122
rect 429 -169 487 -156
rect -487 -338 -429 -325
rect -487 -372 -475 -338
rect -441 -372 -429 -338
rect -487 -406 -429 -372
rect -487 -440 -475 -406
rect -441 -440 -429 -406
rect -487 -474 -429 -440
rect -487 -508 -475 -474
rect -441 -508 -429 -474
rect -487 -542 -429 -508
rect -487 -576 -475 -542
rect -441 -576 -429 -542
rect -487 -610 -429 -576
rect -487 -644 -475 -610
rect -441 -644 -429 -610
rect -487 -678 -429 -644
rect -487 -712 -475 -678
rect -441 -712 -429 -678
rect -487 -725 -429 -712
rect -29 -338 29 -325
rect -29 -372 -17 -338
rect 17 -372 29 -338
rect -29 -406 29 -372
rect -29 -440 -17 -406
rect 17 -440 29 -406
rect -29 -474 29 -440
rect -29 -508 -17 -474
rect 17 -508 29 -474
rect -29 -542 29 -508
rect -29 -576 -17 -542
rect 17 -576 29 -542
rect -29 -610 29 -576
rect -29 -644 -17 -610
rect 17 -644 29 -610
rect -29 -678 29 -644
rect -29 -712 -17 -678
rect 17 -712 29 -678
rect -29 -725 29 -712
rect 429 -338 487 -325
rect 429 -372 441 -338
rect 475 -372 487 -338
rect 429 -406 487 -372
rect 429 -440 441 -406
rect 475 -440 487 -406
rect 429 -474 487 -440
rect 429 -508 441 -474
rect 475 -508 487 -474
rect 429 -542 487 -508
rect 429 -576 441 -542
rect 475 -576 487 -542
rect 429 -610 487 -576
rect 429 -644 441 -610
rect 475 -644 487 -610
rect 429 -678 487 -644
rect 429 -712 441 -678
rect 475 -712 487 -678
rect 429 -725 487 -712
rect -487 -894 -429 -881
rect -487 -928 -475 -894
rect -441 -928 -429 -894
rect -487 -962 -429 -928
rect -487 -996 -475 -962
rect -441 -996 -429 -962
rect -487 -1030 -429 -996
rect -487 -1064 -475 -1030
rect -441 -1064 -429 -1030
rect -487 -1098 -429 -1064
rect -487 -1132 -475 -1098
rect -441 -1132 -429 -1098
rect -487 -1166 -429 -1132
rect -487 -1200 -475 -1166
rect -441 -1200 -429 -1166
rect -487 -1234 -429 -1200
rect -487 -1268 -475 -1234
rect -441 -1268 -429 -1234
rect -487 -1281 -429 -1268
rect -29 -894 29 -881
rect -29 -928 -17 -894
rect 17 -928 29 -894
rect -29 -962 29 -928
rect -29 -996 -17 -962
rect 17 -996 29 -962
rect -29 -1030 29 -996
rect -29 -1064 -17 -1030
rect 17 -1064 29 -1030
rect -29 -1098 29 -1064
rect -29 -1132 -17 -1098
rect 17 -1132 29 -1098
rect -29 -1166 29 -1132
rect -29 -1200 -17 -1166
rect 17 -1200 29 -1166
rect -29 -1234 29 -1200
rect -29 -1268 -17 -1234
rect 17 -1268 29 -1234
rect -29 -1281 29 -1268
rect 429 -894 487 -881
rect 429 -928 441 -894
rect 475 -928 487 -894
rect 429 -962 487 -928
rect 429 -996 441 -962
rect 475 -996 487 -962
rect 429 -1030 487 -996
rect 429 -1064 441 -1030
rect 475 -1064 487 -1030
rect 429 -1098 487 -1064
rect 429 -1132 441 -1098
rect 475 -1132 487 -1098
rect 429 -1166 487 -1132
rect 429 -1200 441 -1166
rect 475 -1200 487 -1166
rect 429 -1234 487 -1200
rect 429 -1268 441 -1234
rect 475 -1268 487 -1234
rect 429 -1281 487 -1268
<< ndiffc >>
rect -475 1296 -441 1330
rect -475 1228 -441 1262
rect -475 1160 -441 1194
rect -475 1092 -441 1126
rect -475 1024 -441 1058
rect -475 956 -441 990
rect -17 1296 17 1330
rect -17 1228 17 1262
rect -17 1160 17 1194
rect -17 1092 17 1126
rect -17 1024 17 1058
rect -17 956 17 990
rect 441 1296 475 1330
rect 441 1228 475 1262
rect 441 1160 475 1194
rect 441 1092 475 1126
rect 441 1024 475 1058
rect 441 956 475 990
rect -475 740 -441 774
rect -475 672 -441 706
rect -475 604 -441 638
rect -475 536 -441 570
rect -475 468 -441 502
rect -475 400 -441 434
rect -17 740 17 774
rect -17 672 17 706
rect -17 604 17 638
rect -17 536 17 570
rect -17 468 17 502
rect -17 400 17 434
rect 441 740 475 774
rect 441 672 475 706
rect 441 604 475 638
rect 441 536 475 570
rect 441 468 475 502
rect 441 400 475 434
rect -475 184 -441 218
rect -475 116 -441 150
rect -475 48 -441 82
rect -475 -20 -441 14
rect -475 -88 -441 -54
rect -475 -156 -441 -122
rect -17 184 17 218
rect -17 116 17 150
rect -17 48 17 82
rect -17 -20 17 14
rect -17 -88 17 -54
rect -17 -156 17 -122
rect 441 184 475 218
rect 441 116 475 150
rect 441 48 475 82
rect 441 -20 475 14
rect 441 -88 475 -54
rect 441 -156 475 -122
rect -475 -372 -441 -338
rect -475 -440 -441 -406
rect -475 -508 -441 -474
rect -475 -576 -441 -542
rect -475 -644 -441 -610
rect -475 -712 -441 -678
rect -17 -372 17 -338
rect -17 -440 17 -406
rect -17 -508 17 -474
rect -17 -576 17 -542
rect -17 -644 17 -610
rect -17 -712 17 -678
rect 441 -372 475 -338
rect 441 -440 475 -406
rect 441 -508 475 -474
rect 441 -576 475 -542
rect 441 -644 475 -610
rect 441 -712 475 -678
rect -475 -928 -441 -894
rect -475 -996 -441 -962
rect -475 -1064 -441 -1030
rect -475 -1132 -441 -1098
rect -475 -1200 -441 -1166
rect -475 -1268 -441 -1234
rect -17 -928 17 -894
rect -17 -996 17 -962
rect -17 -1064 17 -1030
rect -17 -1132 17 -1098
rect -17 -1200 17 -1166
rect -17 -1268 17 -1234
rect 441 -928 475 -894
rect 441 -996 475 -962
rect 441 -1064 475 -1030
rect 441 -1132 475 -1098
rect 441 -1200 475 -1166
rect 441 -1268 475 -1234
<< psubdiff >>
rect -589 1421 -493 1455
rect -459 1421 -425 1455
rect -391 1421 -357 1455
rect -323 1421 -289 1455
rect -255 1421 -221 1455
rect -187 1421 -153 1455
rect -119 1421 -85 1455
rect -51 1421 -17 1455
rect 17 1421 51 1455
rect 85 1421 119 1455
rect 153 1421 187 1455
rect 221 1421 255 1455
rect 289 1421 323 1455
rect 357 1421 391 1455
rect 425 1421 459 1455
rect 493 1421 589 1455
rect -589 1343 -555 1421
rect 555 1343 589 1421
rect -589 1275 -555 1309
rect -589 1207 -555 1241
rect -589 1139 -555 1173
rect -589 1071 -555 1105
rect -589 1003 -555 1037
rect -589 935 -555 969
rect 555 1275 589 1309
rect 555 1207 589 1241
rect 555 1139 589 1173
rect 555 1071 589 1105
rect 555 1003 589 1037
rect -589 867 -555 901
rect 555 935 589 969
rect 555 867 589 901
rect -589 799 -555 833
rect 555 799 589 833
rect -589 731 -555 765
rect -589 663 -555 697
rect -589 595 -555 629
rect -589 527 -555 561
rect -589 459 -555 493
rect -589 391 -555 425
rect 555 731 589 765
rect 555 663 589 697
rect 555 595 589 629
rect 555 527 589 561
rect 555 459 589 493
rect 555 391 589 425
rect -589 323 -555 357
rect 555 323 589 357
rect -589 255 -555 289
rect 555 255 589 289
rect -589 187 -555 221
rect -589 119 -555 153
rect -589 51 -555 85
rect -589 -17 -555 17
rect -589 -85 -555 -51
rect -589 -153 -555 -119
rect 555 187 589 221
rect 555 119 589 153
rect 555 51 589 85
rect 555 -17 589 17
rect 555 -85 589 -51
rect 555 -153 589 -119
rect -589 -221 -555 -187
rect -589 -289 -555 -255
rect 555 -221 589 -187
rect 555 -289 589 -255
rect -589 -357 -555 -323
rect -589 -425 -555 -391
rect -589 -493 -555 -459
rect -589 -561 -555 -527
rect -589 -629 -555 -595
rect -589 -697 -555 -663
rect 555 -357 589 -323
rect 555 -425 589 -391
rect 555 -493 589 -459
rect 555 -561 589 -527
rect 555 -629 589 -595
rect 555 -697 589 -663
rect -589 -765 -555 -731
rect -589 -833 -555 -799
rect 555 -765 589 -731
rect 555 -833 589 -799
rect -589 -901 -555 -867
rect -589 -969 -555 -935
rect -589 -1037 -555 -1003
rect -589 -1105 -555 -1071
rect -589 -1173 -555 -1139
rect -589 -1241 -555 -1207
rect -589 -1309 -555 -1275
rect 555 -901 589 -867
rect 555 -969 589 -935
rect 555 -1037 589 -1003
rect 555 -1105 589 -1071
rect 555 -1173 589 -1139
rect 555 -1241 589 -1207
rect -589 -1421 -555 -1343
rect 555 -1309 589 -1275
rect 555 -1421 589 -1343
rect -589 -1455 -493 -1421
rect -459 -1455 -425 -1421
rect -391 -1455 -357 -1421
rect -323 -1455 -289 -1421
rect -255 -1455 -221 -1421
rect -187 -1455 -153 -1421
rect -119 -1455 -85 -1421
rect -51 -1455 -17 -1421
rect 17 -1455 51 -1421
rect 85 -1455 119 -1421
rect 153 -1455 187 -1421
rect 221 -1455 255 -1421
rect 289 -1455 323 -1421
rect 357 -1455 391 -1421
rect 425 -1455 459 -1421
rect 493 -1455 589 -1421
<< psubdiffcont >>
rect -493 1421 -459 1455
rect -425 1421 -391 1455
rect -357 1421 -323 1455
rect -289 1421 -255 1455
rect -221 1421 -187 1455
rect -153 1421 -119 1455
rect -85 1421 -51 1455
rect -17 1421 17 1455
rect 51 1421 85 1455
rect 119 1421 153 1455
rect 187 1421 221 1455
rect 255 1421 289 1455
rect 323 1421 357 1455
rect 391 1421 425 1455
rect 459 1421 493 1455
rect -589 1309 -555 1343
rect -589 1241 -555 1275
rect -589 1173 -555 1207
rect -589 1105 -555 1139
rect -589 1037 -555 1071
rect -589 969 -555 1003
rect 555 1309 589 1343
rect 555 1241 589 1275
rect 555 1173 589 1207
rect 555 1105 589 1139
rect 555 1037 589 1071
rect 555 969 589 1003
rect -589 901 -555 935
rect -589 833 -555 867
rect 555 901 589 935
rect 555 833 589 867
rect -589 765 -555 799
rect -589 697 -555 731
rect -589 629 -555 663
rect -589 561 -555 595
rect -589 493 -555 527
rect -589 425 -555 459
rect -589 357 -555 391
rect 555 765 589 799
rect 555 697 589 731
rect 555 629 589 663
rect 555 561 589 595
rect 555 493 589 527
rect 555 425 589 459
rect -589 289 -555 323
rect 555 357 589 391
rect 555 289 589 323
rect -589 221 -555 255
rect -589 153 -555 187
rect -589 85 -555 119
rect -589 17 -555 51
rect -589 -51 -555 -17
rect -589 -119 -555 -85
rect -589 -187 -555 -153
rect 555 221 589 255
rect 555 153 589 187
rect 555 85 589 119
rect 555 17 589 51
rect 555 -51 589 -17
rect 555 -119 589 -85
rect -589 -255 -555 -221
rect 555 -187 589 -153
rect 555 -255 589 -221
rect -589 -323 -555 -289
rect 555 -323 589 -289
rect -589 -391 -555 -357
rect -589 -459 -555 -425
rect -589 -527 -555 -493
rect -589 -595 -555 -561
rect -589 -663 -555 -629
rect -589 -731 -555 -697
rect 555 -391 589 -357
rect 555 -459 589 -425
rect 555 -527 589 -493
rect 555 -595 589 -561
rect 555 -663 589 -629
rect -589 -799 -555 -765
rect 555 -731 589 -697
rect 555 -799 589 -765
rect -589 -867 -555 -833
rect 555 -867 589 -833
rect -589 -935 -555 -901
rect -589 -1003 -555 -969
rect -589 -1071 -555 -1037
rect -589 -1139 -555 -1105
rect -589 -1207 -555 -1173
rect -589 -1275 -555 -1241
rect 555 -935 589 -901
rect 555 -1003 589 -969
rect 555 -1071 589 -1037
rect 555 -1139 589 -1105
rect 555 -1207 589 -1173
rect 555 -1275 589 -1241
rect -589 -1343 -555 -1309
rect 555 -1343 589 -1309
rect -493 -1455 -459 -1421
rect -425 -1455 -391 -1421
rect -357 -1455 -323 -1421
rect -289 -1455 -255 -1421
rect -221 -1455 -187 -1421
rect -153 -1455 -119 -1421
rect -85 -1455 -51 -1421
rect -17 -1455 17 -1421
rect 51 -1455 85 -1421
rect 119 -1455 153 -1421
rect 187 -1455 221 -1421
rect 255 -1455 289 -1421
rect 323 -1455 357 -1421
rect 391 -1455 425 -1421
rect 459 -1455 493 -1421
<< poly >>
rect -429 1343 -29 1369
rect 29 1343 429 1369
rect -429 905 -29 943
rect -429 871 -382 905
rect -348 871 -314 905
rect -280 871 -246 905
rect -212 871 -178 905
rect -144 871 -110 905
rect -76 871 -29 905
rect -429 855 -29 871
rect 29 905 429 943
rect 29 871 76 905
rect 110 871 144 905
rect 178 871 212 905
rect 246 871 280 905
rect 314 871 348 905
rect 382 871 429 905
rect 29 855 429 871
rect -429 787 -29 813
rect 29 787 429 813
rect -429 349 -29 387
rect -429 315 -382 349
rect -348 315 -314 349
rect -280 315 -246 349
rect -212 315 -178 349
rect -144 315 -110 349
rect -76 315 -29 349
rect -429 299 -29 315
rect 29 349 429 387
rect 29 315 76 349
rect 110 315 144 349
rect 178 315 212 349
rect 246 315 280 349
rect 314 315 348 349
rect 382 315 429 349
rect 29 299 429 315
rect -429 231 -29 257
rect 29 231 429 257
rect -429 -207 -29 -169
rect -429 -241 -382 -207
rect -348 -241 -314 -207
rect -280 -241 -246 -207
rect -212 -241 -178 -207
rect -144 -241 -110 -207
rect -76 -241 -29 -207
rect -429 -257 -29 -241
rect 29 -207 429 -169
rect 29 -241 76 -207
rect 110 -241 144 -207
rect 178 -241 212 -207
rect 246 -241 280 -207
rect 314 -241 348 -207
rect 382 -241 429 -207
rect 29 -257 429 -241
rect -429 -325 -29 -299
rect 29 -325 429 -299
rect -429 -763 -29 -725
rect -429 -797 -382 -763
rect -348 -797 -314 -763
rect -280 -797 -246 -763
rect -212 -797 -178 -763
rect -144 -797 -110 -763
rect -76 -797 -29 -763
rect -429 -813 -29 -797
rect 29 -763 429 -725
rect 29 -797 76 -763
rect 110 -797 144 -763
rect 178 -797 212 -763
rect 246 -797 280 -763
rect 314 -797 348 -763
rect 382 -797 429 -763
rect 29 -813 429 -797
rect -429 -881 -29 -855
rect 29 -881 429 -855
rect -429 -1319 -29 -1281
rect -429 -1353 -382 -1319
rect -348 -1353 -314 -1319
rect -280 -1353 -246 -1319
rect -212 -1353 -178 -1319
rect -144 -1353 -110 -1319
rect -76 -1353 -29 -1319
rect -429 -1369 -29 -1353
rect 29 -1319 429 -1281
rect 29 -1353 76 -1319
rect 110 -1353 144 -1319
rect 178 -1353 212 -1319
rect 246 -1353 280 -1319
rect 314 -1353 348 -1319
rect 382 -1353 429 -1319
rect 29 -1369 429 -1353
<< polycont >>
rect -382 871 -348 905
rect -314 871 -280 905
rect -246 871 -212 905
rect -178 871 -144 905
rect -110 871 -76 905
rect 76 871 110 905
rect 144 871 178 905
rect 212 871 246 905
rect 280 871 314 905
rect 348 871 382 905
rect -382 315 -348 349
rect -314 315 -280 349
rect -246 315 -212 349
rect -178 315 -144 349
rect -110 315 -76 349
rect 76 315 110 349
rect 144 315 178 349
rect 212 315 246 349
rect 280 315 314 349
rect 348 315 382 349
rect -382 -241 -348 -207
rect -314 -241 -280 -207
rect -246 -241 -212 -207
rect -178 -241 -144 -207
rect -110 -241 -76 -207
rect 76 -241 110 -207
rect 144 -241 178 -207
rect 212 -241 246 -207
rect 280 -241 314 -207
rect 348 -241 382 -207
rect -382 -797 -348 -763
rect -314 -797 -280 -763
rect -246 -797 -212 -763
rect -178 -797 -144 -763
rect -110 -797 -76 -763
rect 76 -797 110 -763
rect 144 -797 178 -763
rect 212 -797 246 -763
rect 280 -797 314 -763
rect 348 -797 382 -763
rect -382 -1353 -348 -1319
rect -314 -1353 -280 -1319
rect -246 -1353 -212 -1319
rect -178 -1353 -144 -1319
rect -110 -1353 -76 -1319
rect 76 -1353 110 -1319
rect 144 -1353 178 -1319
rect 212 -1353 246 -1319
rect 280 -1353 314 -1319
rect 348 -1353 382 -1319
<< locali >>
rect -589 1421 -493 1455
rect -459 1421 -425 1455
rect -391 1421 -357 1455
rect -323 1421 -289 1455
rect -255 1421 -221 1455
rect -187 1421 -153 1455
rect -119 1421 -85 1455
rect -51 1421 -17 1455
rect 17 1421 51 1455
rect 85 1421 119 1455
rect 153 1421 187 1455
rect 221 1421 255 1455
rect 289 1421 323 1455
rect 357 1421 391 1455
rect 425 1421 459 1455
rect 493 1421 589 1455
rect -589 1343 -555 1421
rect -589 1275 -555 1309
rect -589 1207 -555 1241
rect -589 1139 -555 1173
rect -589 1071 -555 1105
rect -589 1003 -555 1037
rect -589 935 -555 969
rect -475 1330 -441 1347
rect -475 1262 -441 1270
rect -475 1194 -441 1198
rect -475 1088 -441 1092
rect -475 1016 -441 1024
rect -475 939 -441 956
rect -17 1330 17 1347
rect -17 1262 17 1270
rect -17 1194 17 1198
rect -17 1088 17 1092
rect -17 1016 17 1024
rect -17 939 17 956
rect 441 1330 475 1347
rect 441 1262 475 1270
rect 441 1194 475 1198
rect 441 1088 475 1092
rect 441 1016 475 1024
rect 441 939 475 956
rect 555 1343 589 1421
rect 555 1275 589 1309
rect 555 1207 589 1241
rect 555 1139 589 1173
rect 555 1071 589 1105
rect 555 1003 589 1037
rect 555 935 589 969
rect -589 867 -555 901
rect -429 871 -390 905
rect -348 871 -318 905
rect -280 871 -246 905
rect -212 871 -178 905
rect -140 871 -110 905
rect -68 871 -29 905
rect 29 871 68 905
rect 110 871 140 905
rect 178 871 212 905
rect 246 871 280 905
rect 318 871 348 905
rect 390 871 429 905
rect -589 799 -555 833
rect 555 867 589 901
rect 555 799 589 833
rect -589 731 -555 765
rect -589 663 -555 697
rect -589 595 -555 629
rect -589 527 -555 561
rect -589 459 -555 493
rect -589 391 -555 425
rect -475 774 -441 791
rect -475 706 -441 714
rect -475 638 -441 642
rect -475 532 -441 536
rect -475 460 -441 468
rect -475 383 -441 400
rect -17 774 17 791
rect -17 706 17 714
rect -17 638 17 642
rect -17 532 17 536
rect -17 460 17 468
rect -17 383 17 400
rect 441 774 475 791
rect 441 706 475 714
rect 441 638 475 642
rect 441 532 475 536
rect 441 460 475 468
rect 441 383 475 400
rect 555 731 589 765
rect 555 663 589 697
rect 555 595 589 629
rect 555 527 589 561
rect 555 459 589 493
rect 555 391 589 425
rect -589 323 -555 357
rect -429 315 -390 349
rect -348 315 -318 349
rect -280 315 -246 349
rect -212 315 -178 349
rect -140 315 -110 349
rect -68 315 -29 349
rect 29 315 68 349
rect 110 315 140 349
rect 178 315 212 349
rect 246 315 280 349
rect 318 315 348 349
rect 390 315 429 349
rect 555 323 589 357
rect -589 255 -555 289
rect 555 255 589 289
rect -589 187 -555 221
rect -589 119 -555 153
rect -589 51 -555 85
rect -589 -17 -555 17
rect -589 -85 -555 -51
rect -589 -153 -555 -119
rect -475 218 -441 235
rect -475 150 -441 158
rect -475 82 -441 86
rect -475 -24 -441 -20
rect -475 -96 -441 -88
rect -475 -173 -441 -156
rect -17 218 17 235
rect -17 150 17 158
rect -17 82 17 86
rect -17 -24 17 -20
rect -17 -96 17 -88
rect -17 -173 17 -156
rect 441 218 475 235
rect 441 150 475 158
rect 441 82 475 86
rect 441 -24 475 -20
rect 441 -96 475 -88
rect 441 -173 475 -156
rect 555 187 589 221
rect 555 119 589 153
rect 555 51 589 85
rect 555 -17 589 17
rect 555 -85 589 -51
rect 555 -153 589 -119
rect -589 -221 -555 -187
rect -429 -241 -390 -207
rect -348 -241 -318 -207
rect -280 -241 -246 -207
rect -212 -241 -178 -207
rect -140 -241 -110 -207
rect -68 -241 -29 -207
rect 29 -241 68 -207
rect 110 -241 140 -207
rect 178 -241 212 -207
rect 246 -241 280 -207
rect 318 -241 348 -207
rect 390 -241 429 -207
rect 555 -221 589 -187
rect -589 -289 -555 -255
rect 555 -289 589 -255
rect -589 -357 -555 -323
rect -589 -425 -555 -391
rect -589 -493 -555 -459
rect -589 -561 -555 -527
rect -589 -629 -555 -595
rect -589 -697 -555 -663
rect -475 -338 -441 -321
rect -475 -406 -441 -398
rect -475 -474 -441 -470
rect -475 -580 -441 -576
rect -475 -652 -441 -644
rect -475 -729 -441 -712
rect -17 -338 17 -321
rect -17 -406 17 -398
rect -17 -474 17 -470
rect -17 -580 17 -576
rect -17 -652 17 -644
rect -17 -729 17 -712
rect 441 -338 475 -321
rect 441 -406 475 -398
rect 441 -474 475 -470
rect 441 -580 475 -576
rect 441 -652 475 -644
rect 441 -729 475 -712
rect 555 -357 589 -323
rect 555 -425 589 -391
rect 555 -493 589 -459
rect 555 -561 589 -527
rect 555 -629 589 -595
rect 555 -697 589 -663
rect -589 -765 -555 -731
rect -429 -797 -390 -763
rect -348 -797 -318 -763
rect -280 -797 -246 -763
rect -212 -797 -178 -763
rect -140 -797 -110 -763
rect -68 -797 -29 -763
rect 29 -797 68 -763
rect 110 -797 140 -763
rect 178 -797 212 -763
rect 246 -797 280 -763
rect 318 -797 348 -763
rect 390 -797 429 -763
rect 555 -765 589 -731
rect -589 -833 -555 -799
rect -589 -901 -555 -867
rect 555 -833 589 -799
rect -589 -969 -555 -935
rect -589 -1037 -555 -1003
rect -589 -1105 -555 -1071
rect -589 -1173 -555 -1139
rect -589 -1241 -555 -1207
rect -589 -1309 -555 -1275
rect -475 -894 -441 -877
rect -475 -962 -441 -954
rect -475 -1030 -441 -1026
rect -475 -1136 -441 -1132
rect -475 -1208 -441 -1200
rect -475 -1285 -441 -1268
rect -17 -894 17 -877
rect -17 -962 17 -954
rect -17 -1030 17 -1026
rect -17 -1136 17 -1132
rect -17 -1208 17 -1200
rect -17 -1285 17 -1268
rect 441 -894 475 -877
rect 441 -962 475 -954
rect 441 -1030 475 -1026
rect 441 -1136 475 -1132
rect 441 -1208 475 -1200
rect 441 -1285 475 -1268
rect 555 -901 589 -867
rect 555 -969 589 -935
rect 555 -1037 589 -1003
rect 555 -1105 589 -1071
rect 555 -1173 589 -1139
rect 555 -1241 589 -1207
rect 555 -1309 589 -1275
rect -589 -1421 -555 -1343
rect -429 -1353 -390 -1319
rect -348 -1353 -318 -1319
rect -280 -1353 -246 -1319
rect -212 -1353 -178 -1319
rect -140 -1353 -110 -1319
rect -68 -1353 -29 -1319
rect 29 -1353 68 -1319
rect 110 -1353 140 -1319
rect 178 -1353 212 -1319
rect 246 -1353 280 -1319
rect 318 -1353 348 -1319
rect 390 -1353 429 -1319
rect 555 -1421 589 -1343
rect -589 -1455 -493 -1421
rect -459 -1455 -425 -1421
rect -391 -1455 -357 -1421
rect -323 -1455 -289 -1421
rect -255 -1455 -221 -1421
rect -187 -1455 -153 -1421
rect -119 -1455 -85 -1421
rect -51 -1455 -17 -1421
rect 17 -1455 51 -1421
rect 85 -1455 119 -1421
rect 153 -1455 187 -1421
rect 221 -1455 255 -1421
rect 289 -1455 323 -1421
rect 357 -1455 391 -1421
rect 425 -1455 459 -1421
rect 493 -1455 589 -1421
<< viali >>
rect -475 1296 -441 1304
rect -475 1270 -441 1296
rect -475 1228 -441 1232
rect -475 1198 -441 1228
rect -475 1126 -441 1160
rect -475 1058 -441 1088
rect -475 1054 -441 1058
rect -475 990 -441 1016
rect -475 982 -441 990
rect -17 1296 17 1304
rect -17 1270 17 1296
rect -17 1228 17 1232
rect -17 1198 17 1228
rect -17 1126 17 1160
rect -17 1058 17 1088
rect -17 1054 17 1058
rect -17 990 17 1016
rect -17 982 17 990
rect 441 1296 475 1304
rect 441 1270 475 1296
rect 441 1228 475 1232
rect 441 1198 475 1228
rect 441 1126 475 1160
rect 441 1058 475 1088
rect 441 1054 475 1058
rect 441 990 475 1016
rect 441 982 475 990
rect -390 871 -382 905
rect -382 871 -356 905
rect -318 871 -314 905
rect -314 871 -284 905
rect -246 871 -212 905
rect -174 871 -144 905
rect -144 871 -140 905
rect -102 871 -76 905
rect -76 871 -68 905
rect 68 871 76 905
rect 76 871 102 905
rect 140 871 144 905
rect 144 871 174 905
rect 212 871 246 905
rect 284 871 314 905
rect 314 871 318 905
rect 356 871 382 905
rect 382 871 390 905
rect -475 740 -441 748
rect -475 714 -441 740
rect -475 672 -441 676
rect -475 642 -441 672
rect -475 570 -441 604
rect -475 502 -441 532
rect -475 498 -441 502
rect -475 434 -441 460
rect -475 426 -441 434
rect -17 740 17 748
rect -17 714 17 740
rect -17 672 17 676
rect -17 642 17 672
rect -17 570 17 604
rect -17 502 17 532
rect -17 498 17 502
rect -17 434 17 460
rect -17 426 17 434
rect 441 740 475 748
rect 441 714 475 740
rect 441 672 475 676
rect 441 642 475 672
rect 441 570 475 604
rect 441 502 475 532
rect 441 498 475 502
rect 441 434 475 460
rect 441 426 475 434
rect -390 315 -382 349
rect -382 315 -356 349
rect -318 315 -314 349
rect -314 315 -284 349
rect -246 315 -212 349
rect -174 315 -144 349
rect -144 315 -140 349
rect -102 315 -76 349
rect -76 315 -68 349
rect 68 315 76 349
rect 76 315 102 349
rect 140 315 144 349
rect 144 315 174 349
rect 212 315 246 349
rect 284 315 314 349
rect 314 315 318 349
rect 356 315 382 349
rect 382 315 390 349
rect -475 184 -441 192
rect -475 158 -441 184
rect -475 116 -441 120
rect -475 86 -441 116
rect -475 14 -441 48
rect -475 -54 -441 -24
rect -475 -58 -441 -54
rect -475 -122 -441 -96
rect -475 -130 -441 -122
rect -17 184 17 192
rect -17 158 17 184
rect -17 116 17 120
rect -17 86 17 116
rect -17 14 17 48
rect -17 -54 17 -24
rect -17 -58 17 -54
rect -17 -122 17 -96
rect -17 -130 17 -122
rect 441 184 475 192
rect 441 158 475 184
rect 441 116 475 120
rect 441 86 475 116
rect 441 14 475 48
rect 441 -54 475 -24
rect 441 -58 475 -54
rect 441 -122 475 -96
rect 441 -130 475 -122
rect -390 -241 -382 -207
rect -382 -241 -356 -207
rect -318 -241 -314 -207
rect -314 -241 -284 -207
rect -246 -241 -212 -207
rect -174 -241 -144 -207
rect -144 -241 -140 -207
rect -102 -241 -76 -207
rect -76 -241 -68 -207
rect 68 -241 76 -207
rect 76 -241 102 -207
rect 140 -241 144 -207
rect 144 -241 174 -207
rect 212 -241 246 -207
rect 284 -241 314 -207
rect 314 -241 318 -207
rect 356 -241 382 -207
rect 382 -241 390 -207
rect -475 -372 -441 -364
rect -475 -398 -441 -372
rect -475 -440 -441 -436
rect -475 -470 -441 -440
rect -475 -542 -441 -508
rect -475 -610 -441 -580
rect -475 -614 -441 -610
rect -475 -678 -441 -652
rect -475 -686 -441 -678
rect -17 -372 17 -364
rect -17 -398 17 -372
rect -17 -440 17 -436
rect -17 -470 17 -440
rect -17 -542 17 -508
rect -17 -610 17 -580
rect -17 -614 17 -610
rect -17 -678 17 -652
rect -17 -686 17 -678
rect 441 -372 475 -364
rect 441 -398 475 -372
rect 441 -440 475 -436
rect 441 -470 475 -440
rect 441 -542 475 -508
rect 441 -610 475 -580
rect 441 -614 475 -610
rect 441 -678 475 -652
rect 441 -686 475 -678
rect -390 -797 -382 -763
rect -382 -797 -356 -763
rect -318 -797 -314 -763
rect -314 -797 -284 -763
rect -246 -797 -212 -763
rect -174 -797 -144 -763
rect -144 -797 -140 -763
rect -102 -797 -76 -763
rect -76 -797 -68 -763
rect 68 -797 76 -763
rect 76 -797 102 -763
rect 140 -797 144 -763
rect 144 -797 174 -763
rect 212 -797 246 -763
rect 284 -797 314 -763
rect 314 -797 318 -763
rect 356 -797 382 -763
rect 382 -797 390 -763
rect -475 -928 -441 -920
rect -475 -954 -441 -928
rect -475 -996 -441 -992
rect -475 -1026 -441 -996
rect -475 -1098 -441 -1064
rect -475 -1166 -441 -1136
rect -475 -1170 -441 -1166
rect -475 -1234 -441 -1208
rect -475 -1242 -441 -1234
rect -17 -928 17 -920
rect -17 -954 17 -928
rect -17 -996 17 -992
rect -17 -1026 17 -996
rect -17 -1098 17 -1064
rect -17 -1166 17 -1136
rect -17 -1170 17 -1166
rect -17 -1234 17 -1208
rect -17 -1242 17 -1234
rect 441 -928 475 -920
rect 441 -954 475 -928
rect 441 -996 475 -992
rect 441 -1026 475 -996
rect 441 -1098 475 -1064
rect 441 -1166 475 -1136
rect 441 -1170 475 -1166
rect 441 -1234 475 -1208
rect 441 -1242 475 -1234
rect -390 -1353 -382 -1319
rect -382 -1353 -356 -1319
rect -318 -1353 -314 -1319
rect -314 -1353 -284 -1319
rect -246 -1353 -212 -1319
rect -174 -1353 -144 -1319
rect -144 -1353 -140 -1319
rect -102 -1353 -76 -1319
rect -76 -1353 -68 -1319
rect 68 -1353 76 -1319
rect 76 -1353 102 -1319
rect 140 -1353 144 -1319
rect 144 -1353 174 -1319
rect 212 -1353 246 -1319
rect 284 -1353 314 -1319
rect 314 -1353 318 -1319
rect 356 -1353 382 -1319
rect 382 -1353 390 -1319
<< metal1 >>
rect -481 1304 -435 1343
rect -481 1270 -475 1304
rect -441 1270 -435 1304
rect -481 1232 -435 1270
rect -481 1198 -475 1232
rect -441 1198 -435 1232
rect -481 1160 -435 1198
rect -481 1126 -475 1160
rect -441 1126 -435 1160
rect -481 1088 -435 1126
rect -481 1054 -475 1088
rect -441 1054 -435 1088
rect -481 1016 -435 1054
rect -481 982 -475 1016
rect -441 982 -435 1016
rect -481 943 -435 982
rect -23 1304 23 1343
rect -23 1270 -17 1304
rect 17 1270 23 1304
rect -23 1232 23 1270
rect -23 1198 -17 1232
rect 17 1198 23 1232
rect -23 1160 23 1198
rect -23 1126 -17 1160
rect 17 1126 23 1160
rect -23 1088 23 1126
rect -23 1054 -17 1088
rect 17 1054 23 1088
rect -23 1016 23 1054
rect -23 982 -17 1016
rect 17 982 23 1016
rect -23 943 23 982
rect 435 1304 481 1343
rect 435 1270 441 1304
rect 475 1270 481 1304
rect 435 1232 481 1270
rect 435 1198 441 1232
rect 475 1198 481 1232
rect 435 1160 481 1198
rect 435 1126 441 1160
rect 475 1126 481 1160
rect 435 1088 481 1126
rect 435 1054 441 1088
rect 475 1054 481 1088
rect 435 1016 481 1054
rect 435 982 441 1016
rect 475 982 481 1016
rect 435 943 481 982
rect -425 905 -33 911
rect -425 871 -390 905
rect -356 871 -318 905
rect -284 871 -246 905
rect -212 871 -174 905
rect -140 871 -102 905
rect -68 871 -33 905
rect -425 865 -33 871
rect 33 905 425 911
rect 33 871 68 905
rect 102 871 140 905
rect 174 871 212 905
rect 246 871 284 905
rect 318 871 356 905
rect 390 871 425 905
rect 33 865 425 871
rect -481 748 -435 787
rect -481 714 -475 748
rect -441 714 -435 748
rect -481 676 -435 714
rect -481 642 -475 676
rect -441 642 -435 676
rect -481 604 -435 642
rect -481 570 -475 604
rect -441 570 -435 604
rect -481 532 -435 570
rect -481 498 -475 532
rect -441 498 -435 532
rect -481 460 -435 498
rect -481 426 -475 460
rect -441 426 -435 460
rect -481 387 -435 426
rect -23 748 23 787
rect -23 714 -17 748
rect 17 714 23 748
rect -23 676 23 714
rect -23 642 -17 676
rect 17 642 23 676
rect -23 604 23 642
rect -23 570 -17 604
rect 17 570 23 604
rect -23 532 23 570
rect -23 498 -17 532
rect 17 498 23 532
rect -23 460 23 498
rect -23 426 -17 460
rect 17 426 23 460
rect -23 387 23 426
rect 435 748 481 787
rect 435 714 441 748
rect 475 714 481 748
rect 435 676 481 714
rect 435 642 441 676
rect 475 642 481 676
rect 435 604 481 642
rect 435 570 441 604
rect 475 570 481 604
rect 435 532 481 570
rect 435 498 441 532
rect 475 498 481 532
rect 435 460 481 498
rect 435 426 441 460
rect 475 426 481 460
rect 435 387 481 426
rect -425 349 -33 355
rect -425 315 -390 349
rect -356 315 -318 349
rect -284 315 -246 349
rect -212 315 -174 349
rect -140 315 -102 349
rect -68 315 -33 349
rect -425 309 -33 315
rect 33 349 425 355
rect 33 315 68 349
rect 102 315 140 349
rect 174 315 212 349
rect 246 315 284 349
rect 318 315 356 349
rect 390 315 425 349
rect 33 309 425 315
rect -481 192 -435 231
rect -481 158 -475 192
rect -441 158 -435 192
rect -481 120 -435 158
rect -481 86 -475 120
rect -441 86 -435 120
rect -481 48 -435 86
rect -481 14 -475 48
rect -441 14 -435 48
rect -481 -24 -435 14
rect -481 -58 -475 -24
rect -441 -58 -435 -24
rect -481 -96 -435 -58
rect -481 -130 -475 -96
rect -441 -130 -435 -96
rect -481 -169 -435 -130
rect -23 192 23 231
rect -23 158 -17 192
rect 17 158 23 192
rect -23 120 23 158
rect -23 86 -17 120
rect 17 86 23 120
rect -23 48 23 86
rect -23 14 -17 48
rect 17 14 23 48
rect -23 -24 23 14
rect -23 -58 -17 -24
rect 17 -58 23 -24
rect -23 -96 23 -58
rect -23 -130 -17 -96
rect 17 -130 23 -96
rect -23 -169 23 -130
rect 435 192 481 231
rect 435 158 441 192
rect 475 158 481 192
rect 435 120 481 158
rect 435 86 441 120
rect 475 86 481 120
rect 435 48 481 86
rect 435 14 441 48
rect 475 14 481 48
rect 435 -24 481 14
rect 435 -58 441 -24
rect 475 -58 481 -24
rect 435 -96 481 -58
rect 435 -130 441 -96
rect 475 -130 481 -96
rect 435 -169 481 -130
rect -425 -207 -33 -201
rect -425 -241 -390 -207
rect -356 -241 -318 -207
rect -284 -241 -246 -207
rect -212 -241 -174 -207
rect -140 -241 -102 -207
rect -68 -241 -33 -207
rect -425 -247 -33 -241
rect 33 -207 425 -201
rect 33 -241 68 -207
rect 102 -241 140 -207
rect 174 -241 212 -207
rect 246 -241 284 -207
rect 318 -241 356 -207
rect 390 -241 425 -207
rect 33 -247 425 -241
rect -481 -364 -435 -325
rect -481 -398 -475 -364
rect -441 -398 -435 -364
rect -481 -436 -435 -398
rect -481 -470 -475 -436
rect -441 -470 -435 -436
rect -481 -508 -435 -470
rect -481 -542 -475 -508
rect -441 -542 -435 -508
rect -481 -580 -435 -542
rect -481 -614 -475 -580
rect -441 -614 -435 -580
rect -481 -652 -435 -614
rect -481 -686 -475 -652
rect -441 -686 -435 -652
rect -481 -725 -435 -686
rect -23 -364 23 -325
rect -23 -398 -17 -364
rect 17 -398 23 -364
rect -23 -436 23 -398
rect -23 -470 -17 -436
rect 17 -470 23 -436
rect -23 -508 23 -470
rect -23 -542 -17 -508
rect 17 -542 23 -508
rect -23 -580 23 -542
rect -23 -614 -17 -580
rect 17 -614 23 -580
rect -23 -652 23 -614
rect -23 -686 -17 -652
rect 17 -686 23 -652
rect -23 -725 23 -686
rect 435 -364 481 -325
rect 435 -398 441 -364
rect 475 -398 481 -364
rect 435 -436 481 -398
rect 435 -470 441 -436
rect 475 -470 481 -436
rect 435 -508 481 -470
rect 435 -542 441 -508
rect 475 -542 481 -508
rect 435 -580 481 -542
rect 435 -614 441 -580
rect 475 -614 481 -580
rect 435 -652 481 -614
rect 435 -686 441 -652
rect 475 -686 481 -652
rect 435 -725 481 -686
rect -425 -763 -33 -757
rect -425 -797 -390 -763
rect -356 -797 -318 -763
rect -284 -797 -246 -763
rect -212 -797 -174 -763
rect -140 -797 -102 -763
rect -68 -797 -33 -763
rect -425 -803 -33 -797
rect 33 -763 425 -757
rect 33 -797 68 -763
rect 102 -797 140 -763
rect 174 -797 212 -763
rect 246 -797 284 -763
rect 318 -797 356 -763
rect 390 -797 425 -763
rect 33 -803 425 -797
rect -481 -920 -435 -881
rect -481 -954 -475 -920
rect -441 -954 -435 -920
rect -481 -992 -435 -954
rect -481 -1026 -475 -992
rect -441 -1026 -435 -992
rect -481 -1064 -435 -1026
rect -481 -1098 -475 -1064
rect -441 -1098 -435 -1064
rect -481 -1136 -435 -1098
rect -481 -1170 -475 -1136
rect -441 -1170 -435 -1136
rect -481 -1208 -435 -1170
rect -481 -1242 -475 -1208
rect -441 -1242 -435 -1208
rect -481 -1281 -435 -1242
rect -23 -920 23 -881
rect -23 -954 -17 -920
rect 17 -954 23 -920
rect -23 -992 23 -954
rect -23 -1026 -17 -992
rect 17 -1026 23 -992
rect -23 -1064 23 -1026
rect -23 -1098 -17 -1064
rect 17 -1098 23 -1064
rect -23 -1136 23 -1098
rect -23 -1170 -17 -1136
rect 17 -1170 23 -1136
rect -23 -1208 23 -1170
rect -23 -1242 -17 -1208
rect 17 -1242 23 -1208
rect -23 -1281 23 -1242
rect 435 -920 481 -881
rect 435 -954 441 -920
rect 475 -954 481 -920
rect 435 -992 481 -954
rect 435 -1026 441 -992
rect 475 -1026 481 -992
rect 435 -1064 481 -1026
rect 435 -1098 441 -1064
rect 475 -1098 481 -1064
rect 435 -1136 481 -1098
rect 435 -1170 441 -1136
rect 475 -1170 481 -1136
rect 435 -1208 481 -1170
rect 435 -1242 441 -1208
rect 475 -1242 481 -1208
rect 435 -1281 481 -1242
rect -425 -1319 -33 -1313
rect -425 -1353 -390 -1319
rect -356 -1353 -318 -1319
rect -284 -1353 -246 -1319
rect -212 -1353 -174 -1319
rect -140 -1353 -102 -1319
rect -68 -1353 -33 -1319
rect -425 -1359 -33 -1353
rect 33 -1319 425 -1313
rect 33 -1353 68 -1319
rect 102 -1353 140 -1319
rect 174 -1353 212 -1319
rect 246 -1353 284 -1319
rect 318 -1353 356 -1319
rect 390 -1353 425 -1319
rect 33 -1359 425 -1353
<< properties >>
string FIXED_BBOX -572 -1438 572 1438
<< end >>
