magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -968 383 968 634
rect -968 18 968 269
rect -968 -347 968 -96
<< nwell >>
rect -968 383 968 745
rect -968 18 968 380
rect -968 -347 968 15
rect -968 -712 968 -350
<< pmoslvt >>
rect -874 483 -674 683
rect -616 483 -416 683
rect -358 483 -158 683
rect -100 483 100 683
rect 158 483 358 683
rect 416 483 616 683
rect 674 483 874 683
rect -874 118 -674 318
rect -616 118 -416 318
rect -358 118 -158 318
rect -100 118 100 318
rect 158 118 358 318
rect 416 118 616 318
rect 674 118 874 318
rect -874 -247 -674 -47
rect -616 -247 -416 -47
rect -358 -247 -158 -47
rect -100 -247 100 -47
rect 158 -247 358 -47
rect 416 -247 616 -47
rect 674 -247 874 -47
rect -874 -612 -674 -412
rect -616 -612 -416 -412
rect -358 -612 -158 -412
rect -100 -612 100 -412
rect 158 -612 358 -412
rect 416 -612 616 -412
rect 674 -612 874 -412
<< pdiff >>
rect -932 668 -874 683
rect -932 634 -920 668
rect -886 634 -874 668
rect -932 600 -874 634
rect -932 566 -920 600
rect -886 566 -874 600
rect -932 532 -874 566
rect -932 498 -920 532
rect -886 498 -874 532
rect -932 483 -874 498
rect -674 668 -616 683
rect -674 634 -662 668
rect -628 634 -616 668
rect -674 600 -616 634
rect -674 566 -662 600
rect -628 566 -616 600
rect -674 532 -616 566
rect -674 498 -662 532
rect -628 498 -616 532
rect -674 483 -616 498
rect -416 668 -358 683
rect -416 634 -404 668
rect -370 634 -358 668
rect -416 600 -358 634
rect -416 566 -404 600
rect -370 566 -358 600
rect -416 532 -358 566
rect -416 498 -404 532
rect -370 498 -358 532
rect -416 483 -358 498
rect -158 668 -100 683
rect -158 634 -146 668
rect -112 634 -100 668
rect -158 600 -100 634
rect -158 566 -146 600
rect -112 566 -100 600
rect -158 532 -100 566
rect -158 498 -146 532
rect -112 498 -100 532
rect -158 483 -100 498
rect 100 668 158 683
rect 100 634 112 668
rect 146 634 158 668
rect 100 600 158 634
rect 100 566 112 600
rect 146 566 158 600
rect 100 532 158 566
rect 100 498 112 532
rect 146 498 158 532
rect 100 483 158 498
rect 358 668 416 683
rect 358 634 370 668
rect 404 634 416 668
rect 358 600 416 634
rect 358 566 370 600
rect 404 566 416 600
rect 358 532 416 566
rect 358 498 370 532
rect 404 498 416 532
rect 358 483 416 498
rect 616 668 674 683
rect 616 634 628 668
rect 662 634 674 668
rect 616 600 674 634
rect 616 566 628 600
rect 662 566 674 600
rect 616 532 674 566
rect 616 498 628 532
rect 662 498 674 532
rect 616 483 674 498
rect 874 668 932 683
rect 874 634 886 668
rect 920 634 932 668
rect 874 600 932 634
rect 874 566 886 600
rect 920 566 932 600
rect 874 532 932 566
rect 874 498 886 532
rect 920 498 932 532
rect 874 483 932 498
rect -932 303 -874 318
rect -932 269 -920 303
rect -886 269 -874 303
rect -932 235 -874 269
rect -932 201 -920 235
rect -886 201 -874 235
rect -932 167 -874 201
rect -932 133 -920 167
rect -886 133 -874 167
rect -932 118 -874 133
rect -674 303 -616 318
rect -674 269 -662 303
rect -628 269 -616 303
rect -674 235 -616 269
rect -674 201 -662 235
rect -628 201 -616 235
rect -674 167 -616 201
rect -674 133 -662 167
rect -628 133 -616 167
rect -674 118 -616 133
rect -416 303 -358 318
rect -416 269 -404 303
rect -370 269 -358 303
rect -416 235 -358 269
rect -416 201 -404 235
rect -370 201 -358 235
rect -416 167 -358 201
rect -416 133 -404 167
rect -370 133 -358 167
rect -416 118 -358 133
rect -158 303 -100 318
rect -158 269 -146 303
rect -112 269 -100 303
rect -158 235 -100 269
rect -158 201 -146 235
rect -112 201 -100 235
rect -158 167 -100 201
rect -158 133 -146 167
rect -112 133 -100 167
rect -158 118 -100 133
rect 100 303 158 318
rect 100 269 112 303
rect 146 269 158 303
rect 100 235 158 269
rect 100 201 112 235
rect 146 201 158 235
rect 100 167 158 201
rect 100 133 112 167
rect 146 133 158 167
rect 100 118 158 133
rect 358 303 416 318
rect 358 269 370 303
rect 404 269 416 303
rect 358 235 416 269
rect 358 201 370 235
rect 404 201 416 235
rect 358 167 416 201
rect 358 133 370 167
rect 404 133 416 167
rect 358 118 416 133
rect 616 303 674 318
rect 616 269 628 303
rect 662 269 674 303
rect 616 235 674 269
rect 616 201 628 235
rect 662 201 674 235
rect 616 167 674 201
rect 616 133 628 167
rect 662 133 674 167
rect 616 118 674 133
rect 874 303 932 318
rect 874 269 886 303
rect 920 269 932 303
rect 874 235 932 269
rect 874 201 886 235
rect 920 201 932 235
rect 874 167 932 201
rect 874 133 886 167
rect 920 133 932 167
rect 874 118 932 133
rect -932 -62 -874 -47
rect -932 -96 -920 -62
rect -886 -96 -874 -62
rect -932 -130 -874 -96
rect -932 -164 -920 -130
rect -886 -164 -874 -130
rect -932 -198 -874 -164
rect -932 -232 -920 -198
rect -886 -232 -874 -198
rect -932 -247 -874 -232
rect -674 -62 -616 -47
rect -674 -96 -662 -62
rect -628 -96 -616 -62
rect -674 -130 -616 -96
rect -674 -164 -662 -130
rect -628 -164 -616 -130
rect -674 -198 -616 -164
rect -674 -232 -662 -198
rect -628 -232 -616 -198
rect -674 -247 -616 -232
rect -416 -62 -358 -47
rect -416 -96 -404 -62
rect -370 -96 -358 -62
rect -416 -130 -358 -96
rect -416 -164 -404 -130
rect -370 -164 -358 -130
rect -416 -198 -358 -164
rect -416 -232 -404 -198
rect -370 -232 -358 -198
rect -416 -247 -358 -232
rect -158 -62 -100 -47
rect -158 -96 -146 -62
rect -112 -96 -100 -62
rect -158 -130 -100 -96
rect -158 -164 -146 -130
rect -112 -164 -100 -130
rect -158 -198 -100 -164
rect -158 -232 -146 -198
rect -112 -232 -100 -198
rect -158 -247 -100 -232
rect 100 -62 158 -47
rect 100 -96 112 -62
rect 146 -96 158 -62
rect 100 -130 158 -96
rect 100 -164 112 -130
rect 146 -164 158 -130
rect 100 -198 158 -164
rect 100 -232 112 -198
rect 146 -232 158 -198
rect 100 -247 158 -232
rect 358 -62 416 -47
rect 358 -96 370 -62
rect 404 -96 416 -62
rect 358 -130 416 -96
rect 358 -164 370 -130
rect 404 -164 416 -130
rect 358 -198 416 -164
rect 358 -232 370 -198
rect 404 -232 416 -198
rect 358 -247 416 -232
rect 616 -62 674 -47
rect 616 -96 628 -62
rect 662 -96 674 -62
rect 616 -130 674 -96
rect 616 -164 628 -130
rect 662 -164 674 -130
rect 616 -198 674 -164
rect 616 -232 628 -198
rect 662 -232 674 -198
rect 616 -247 674 -232
rect 874 -62 932 -47
rect 874 -96 886 -62
rect 920 -96 932 -62
rect 874 -130 932 -96
rect 874 -164 886 -130
rect 920 -164 932 -130
rect 874 -198 932 -164
rect 874 -232 886 -198
rect 920 -232 932 -198
rect 874 -247 932 -232
rect -932 -427 -874 -412
rect -932 -461 -920 -427
rect -886 -461 -874 -427
rect -932 -495 -874 -461
rect -932 -529 -920 -495
rect -886 -529 -874 -495
rect -932 -563 -874 -529
rect -932 -597 -920 -563
rect -886 -597 -874 -563
rect -932 -612 -874 -597
rect -674 -427 -616 -412
rect -674 -461 -662 -427
rect -628 -461 -616 -427
rect -674 -495 -616 -461
rect -674 -529 -662 -495
rect -628 -529 -616 -495
rect -674 -563 -616 -529
rect -674 -597 -662 -563
rect -628 -597 -616 -563
rect -674 -612 -616 -597
rect -416 -427 -358 -412
rect -416 -461 -404 -427
rect -370 -461 -358 -427
rect -416 -495 -358 -461
rect -416 -529 -404 -495
rect -370 -529 -358 -495
rect -416 -563 -358 -529
rect -416 -597 -404 -563
rect -370 -597 -358 -563
rect -416 -612 -358 -597
rect -158 -427 -100 -412
rect -158 -461 -146 -427
rect -112 -461 -100 -427
rect -158 -495 -100 -461
rect -158 -529 -146 -495
rect -112 -529 -100 -495
rect -158 -563 -100 -529
rect -158 -597 -146 -563
rect -112 -597 -100 -563
rect -158 -612 -100 -597
rect 100 -427 158 -412
rect 100 -461 112 -427
rect 146 -461 158 -427
rect 100 -495 158 -461
rect 100 -529 112 -495
rect 146 -529 158 -495
rect 100 -563 158 -529
rect 100 -597 112 -563
rect 146 -597 158 -563
rect 100 -612 158 -597
rect 358 -427 416 -412
rect 358 -461 370 -427
rect 404 -461 416 -427
rect 358 -495 416 -461
rect 358 -529 370 -495
rect 404 -529 416 -495
rect 358 -563 416 -529
rect 358 -597 370 -563
rect 404 -597 416 -563
rect 358 -612 416 -597
rect 616 -427 674 -412
rect 616 -461 628 -427
rect 662 -461 674 -427
rect 616 -495 674 -461
rect 616 -529 628 -495
rect 662 -529 674 -495
rect 616 -563 674 -529
rect 616 -597 628 -563
rect 662 -597 674 -563
rect 616 -612 674 -597
rect 874 -427 932 -412
rect 874 -461 886 -427
rect 920 -461 932 -427
rect 874 -495 932 -461
rect 874 -529 886 -495
rect 920 -529 932 -495
rect 874 -563 932 -529
rect 874 -597 886 -563
rect 920 -597 932 -563
rect 874 -612 932 -597
<< pdiffc >>
rect -920 634 -886 668
rect -920 566 -886 600
rect -920 498 -886 532
rect -662 634 -628 668
rect -662 566 -628 600
rect -662 498 -628 532
rect -404 634 -370 668
rect -404 566 -370 600
rect -404 498 -370 532
rect -146 634 -112 668
rect -146 566 -112 600
rect -146 498 -112 532
rect 112 634 146 668
rect 112 566 146 600
rect 112 498 146 532
rect 370 634 404 668
rect 370 566 404 600
rect 370 498 404 532
rect 628 634 662 668
rect 628 566 662 600
rect 628 498 662 532
rect 886 634 920 668
rect 886 566 920 600
rect 886 498 920 532
rect -920 269 -886 303
rect -920 201 -886 235
rect -920 133 -886 167
rect -662 269 -628 303
rect -662 201 -628 235
rect -662 133 -628 167
rect -404 269 -370 303
rect -404 201 -370 235
rect -404 133 -370 167
rect -146 269 -112 303
rect -146 201 -112 235
rect -146 133 -112 167
rect 112 269 146 303
rect 112 201 146 235
rect 112 133 146 167
rect 370 269 404 303
rect 370 201 404 235
rect 370 133 404 167
rect 628 269 662 303
rect 628 201 662 235
rect 628 133 662 167
rect 886 269 920 303
rect 886 201 920 235
rect 886 133 920 167
rect -920 -96 -886 -62
rect -920 -164 -886 -130
rect -920 -232 -886 -198
rect -662 -96 -628 -62
rect -662 -164 -628 -130
rect -662 -232 -628 -198
rect -404 -96 -370 -62
rect -404 -164 -370 -130
rect -404 -232 -370 -198
rect -146 -96 -112 -62
rect -146 -164 -112 -130
rect -146 -232 -112 -198
rect 112 -96 146 -62
rect 112 -164 146 -130
rect 112 -232 146 -198
rect 370 -96 404 -62
rect 370 -164 404 -130
rect 370 -232 404 -198
rect 628 -96 662 -62
rect 628 -164 662 -130
rect 628 -232 662 -198
rect 886 -96 920 -62
rect 886 -164 920 -130
rect 886 -232 920 -198
rect -920 -461 -886 -427
rect -920 -529 -886 -495
rect -920 -597 -886 -563
rect -662 -461 -628 -427
rect -662 -529 -628 -495
rect -662 -597 -628 -563
rect -404 -461 -370 -427
rect -404 -529 -370 -495
rect -404 -597 -370 -563
rect -146 -461 -112 -427
rect -146 -529 -112 -495
rect -146 -597 -112 -563
rect 112 -461 146 -427
rect 112 -529 146 -495
rect 112 -597 146 -563
rect 370 -461 404 -427
rect 370 -529 404 -495
rect 370 -597 404 -563
rect 628 -461 662 -427
rect 628 -529 662 -495
rect 628 -597 662 -563
rect 886 -461 920 -427
rect 886 -529 920 -495
rect 886 -597 920 -563
<< poly >>
rect -874 683 -674 709
rect -616 683 -416 709
rect -358 683 -158 709
rect -100 683 100 709
rect 158 683 358 709
rect 416 683 616 709
rect 674 683 874 709
rect -874 436 -674 483
rect -874 402 -825 436
rect -791 402 -757 436
rect -723 402 -674 436
rect -874 386 -674 402
rect -616 436 -416 483
rect -616 402 -567 436
rect -533 402 -499 436
rect -465 402 -416 436
rect -616 386 -416 402
rect -358 436 -158 483
rect -358 402 -309 436
rect -275 402 -241 436
rect -207 402 -158 436
rect -358 386 -158 402
rect -100 436 100 483
rect -100 402 -51 436
rect -17 402 17 436
rect 51 402 100 436
rect -100 386 100 402
rect 158 436 358 483
rect 158 402 207 436
rect 241 402 275 436
rect 309 402 358 436
rect 158 386 358 402
rect 416 436 616 483
rect 416 402 465 436
rect 499 402 533 436
rect 567 402 616 436
rect 416 386 616 402
rect 674 436 874 483
rect 674 402 723 436
rect 757 402 791 436
rect 825 402 874 436
rect 674 386 874 402
rect -874 318 -674 344
rect -616 318 -416 344
rect -358 318 -158 344
rect -100 318 100 344
rect 158 318 358 344
rect 416 318 616 344
rect 674 318 874 344
rect -874 71 -674 118
rect -874 37 -825 71
rect -791 37 -757 71
rect -723 37 -674 71
rect -874 21 -674 37
rect -616 71 -416 118
rect -616 37 -567 71
rect -533 37 -499 71
rect -465 37 -416 71
rect -616 21 -416 37
rect -358 71 -158 118
rect -358 37 -309 71
rect -275 37 -241 71
rect -207 37 -158 71
rect -358 21 -158 37
rect -100 71 100 118
rect -100 37 -51 71
rect -17 37 17 71
rect 51 37 100 71
rect -100 21 100 37
rect 158 71 358 118
rect 158 37 207 71
rect 241 37 275 71
rect 309 37 358 71
rect 158 21 358 37
rect 416 71 616 118
rect 416 37 465 71
rect 499 37 533 71
rect 567 37 616 71
rect 416 21 616 37
rect 674 71 874 118
rect 674 37 723 71
rect 757 37 791 71
rect 825 37 874 71
rect 674 21 874 37
rect -874 -47 -674 -21
rect -616 -47 -416 -21
rect -358 -47 -158 -21
rect -100 -47 100 -21
rect 158 -47 358 -21
rect 416 -47 616 -21
rect 674 -47 874 -21
rect -874 -294 -674 -247
rect -874 -328 -825 -294
rect -791 -328 -757 -294
rect -723 -328 -674 -294
rect -874 -344 -674 -328
rect -616 -294 -416 -247
rect -616 -328 -567 -294
rect -533 -328 -499 -294
rect -465 -328 -416 -294
rect -616 -344 -416 -328
rect -358 -294 -158 -247
rect -358 -328 -309 -294
rect -275 -328 -241 -294
rect -207 -328 -158 -294
rect -358 -344 -158 -328
rect -100 -294 100 -247
rect -100 -328 -51 -294
rect -17 -328 17 -294
rect 51 -328 100 -294
rect -100 -344 100 -328
rect 158 -294 358 -247
rect 158 -328 207 -294
rect 241 -328 275 -294
rect 309 -328 358 -294
rect 158 -344 358 -328
rect 416 -294 616 -247
rect 416 -328 465 -294
rect 499 -328 533 -294
rect 567 -328 616 -294
rect 416 -344 616 -328
rect 674 -294 874 -247
rect 674 -328 723 -294
rect 757 -328 791 -294
rect 825 -328 874 -294
rect 674 -344 874 -328
rect -874 -412 -674 -386
rect -616 -412 -416 -386
rect -358 -412 -158 -386
rect -100 -412 100 -386
rect 158 -412 358 -386
rect 416 -412 616 -386
rect 674 -412 874 -386
rect -874 -659 -674 -612
rect -874 -693 -825 -659
rect -791 -693 -757 -659
rect -723 -693 -674 -659
rect -874 -709 -674 -693
rect -616 -659 -416 -612
rect -616 -693 -567 -659
rect -533 -693 -499 -659
rect -465 -693 -416 -659
rect -616 -709 -416 -693
rect -358 -659 -158 -612
rect -358 -693 -309 -659
rect -275 -693 -241 -659
rect -207 -693 -158 -659
rect -358 -709 -158 -693
rect -100 -659 100 -612
rect -100 -693 -51 -659
rect -17 -693 17 -659
rect 51 -693 100 -659
rect -100 -709 100 -693
rect 158 -659 358 -612
rect 158 -693 207 -659
rect 241 -693 275 -659
rect 309 -693 358 -659
rect 158 -709 358 -693
rect 416 -659 616 -612
rect 416 -693 465 -659
rect 499 -693 533 -659
rect 567 -693 616 -659
rect 416 -709 616 -693
rect 674 -659 874 -612
rect 674 -693 723 -659
rect 757 -693 791 -659
rect 825 -693 874 -659
rect 674 -709 874 -693
<< polycont >>
rect -825 402 -791 436
rect -757 402 -723 436
rect -567 402 -533 436
rect -499 402 -465 436
rect -309 402 -275 436
rect -241 402 -207 436
rect -51 402 -17 436
rect 17 402 51 436
rect 207 402 241 436
rect 275 402 309 436
rect 465 402 499 436
rect 533 402 567 436
rect 723 402 757 436
rect 791 402 825 436
rect -825 37 -791 71
rect -757 37 -723 71
rect -567 37 -533 71
rect -499 37 -465 71
rect -309 37 -275 71
rect -241 37 -207 71
rect -51 37 -17 71
rect 17 37 51 71
rect 207 37 241 71
rect 275 37 309 71
rect 465 37 499 71
rect 533 37 567 71
rect 723 37 757 71
rect 791 37 825 71
rect -825 -328 -791 -294
rect -757 -328 -723 -294
rect -567 -328 -533 -294
rect -499 -328 -465 -294
rect -309 -328 -275 -294
rect -241 -328 -207 -294
rect -51 -328 -17 -294
rect 17 -328 51 -294
rect 207 -328 241 -294
rect 275 -328 309 -294
rect 465 -328 499 -294
rect 533 -328 567 -294
rect 723 -328 757 -294
rect 791 -328 825 -294
rect -825 -693 -791 -659
rect -757 -693 -723 -659
rect -567 -693 -533 -659
rect -499 -693 -465 -659
rect -309 -693 -275 -659
rect -241 -693 -207 -659
rect -51 -693 -17 -659
rect 17 -693 51 -659
rect 207 -693 241 -659
rect 275 -693 309 -659
rect 465 -693 499 -659
rect 533 -693 567 -659
rect 723 -693 757 -659
rect 791 -693 825 -659
<< locali >>
rect -920 668 -886 687
rect -920 600 -886 602
rect -920 564 -886 566
rect -920 479 -886 498
rect -662 668 -628 687
rect -662 600 -628 602
rect -662 564 -628 566
rect -662 479 -628 498
rect -404 668 -370 687
rect -404 600 -370 602
rect -404 564 -370 566
rect -404 479 -370 498
rect -146 668 -112 687
rect -146 600 -112 602
rect -146 564 -112 566
rect -146 479 -112 498
rect 112 668 146 687
rect 112 600 146 602
rect 112 564 146 566
rect 112 479 146 498
rect 370 668 404 687
rect 370 600 404 602
rect 370 564 404 566
rect 370 479 404 498
rect 628 668 662 687
rect 628 600 662 602
rect 628 564 662 566
rect 628 479 662 498
rect 886 668 920 687
rect 886 600 920 602
rect 886 564 920 566
rect 886 479 920 498
rect -874 402 -827 436
rect -791 402 -757 436
rect -721 402 -674 436
rect -616 402 -569 436
rect -533 402 -499 436
rect -463 402 -416 436
rect -358 402 -311 436
rect -275 402 -241 436
rect -205 402 -158 436
rect -100 402 -53 436
rect -17 402 17 436
rect 53 402 100 436
rect 158 402 205 436
rect 241 402 275 436
rect 311 402 358 436
rect 416 402 463 436
rect 499 402 533 436
rect 569 402 616 436
rect 674 402 721 436
rect 757 402 791 436
rect 827 402 874 436
rect -920 303 -886 322
rect -920 235 -886 237
rect -920 199 -886 201
rect -920 114 -886 133
rect -662 303 -628 322
rect -662 235 -628 237
rect -662 199 -628 201
rect -662 114 -628 133
rect -404 303 -370 322
rect -404 235 -370 237
rect -404 199 -370 201
rect -404 114 -370 133
rect -146 303 -112 322
rect -146 235 -112 237
rect -146 199 -112 201
rect -146 114 -112 133
rect 112 303 146 322
rect 112 235 146 237
rect 112 199 146 201
rect 112 114 146 133
rect 370 303 404 322
rect 370 235 404 237
rect 370 199 404 201
rect 370 114 404 133
rect 628 303 662 322
rect 628 235 662 237
rect 628 199 662 201
rect 628 114 662 133
rect 886 303 920 322
rect 886 235 920 237
rect 886 199 920 201
rect 886 114 920 133
rect -874 37 -827 71
rect -791 37 -757 71
rect -721 37 -674 71
rect -616 37 -569 71
rect -533 37 -499 71
rect -463 37 -416 71
rect -358 37 -311 71
rect -275 37 -241 71
rect -205 37 -158 71
rect -100 37 -53 71
rect -17 37 17 71
rect 53 37 100 71
rect 158 37 205 71
rect 241 37 275 71
rect 311 37 358 71
rect 416 37 463 71
rect 499 37 533 71
rect 569 37 616 71
rect 674 37 721 71
rect 757 37 791 71
rect 827 37 874 71
rect -920 -62 -886 -43
rect -920 -130 -886 -128
rect -920 -166 -886 -164
rect -920 -251 -886 -232
rect -662 -62 -628 -43
rect -662 -130 -628 -128
rect -662 -166 -628 -164
rect -662 -251 -628 -232
rect -404 -62 -370 -43
rect -404 -130 -370 -128
rect -404 -166 -370 -164
rect -404 -251 -370 -232
rect -146 -62 -112 -43
rect -146 -130 -112 -128
rect -146 -166 -112 -164
rect -146 -251 -112 -232
rect 112 -62 146 -43
rect 112 -130 146 -128
rect 112 -166 146 -164
rect 112 -251 146 -232
rect 370 -62 404 -43
rect 370 -130 404 -128
rect 370 -166 404 -164
rect 370 -251 404 -232
rect 628 -62 662 -43
rect 628 -130 662 -128
rect 628 -166 662 -164
rect 628 -251 662 -232
rect 886 -62 920 -43
rect 886 -130 920 -128
rect 886 -166 920 -164
rect 886 -251 920 -232
rect -874 -328 -827 -294
rect -791 -328 -757 -294
rect -721 -328 -674 -294
rect -616 -328 -569 -294
rect -533 -328 -499 -294
rect -463 -328 -416 -294
rect -358 -328 -311 -294
rect -275 -328 -241 -294
rect -205 -328 -158 -294
rect -100 -328 -53 -294
rect -17 -328 17 -294
rect 53 -328 100 -294
rect 158 -328 205 -294
rect 241 -328 275 -294
rect 311 -328 358 -294
rect 416 -328 463 -294
rect 499 -328 533 -294
rect 569 -328 616 -294
rect 674 -328 721 -294
rect 757 -328 791 -294
rect 827 -328 874 -294
rect -920 -427 -886 -408
rect -920 -495 -886 -493
rect -920 -531 -886 -529
rect -920 -616 -886 -597
rect -662 -427 -628 -408
rect -662 -495 -628 -493
rect -662 -531 -628 -529
rect -662 -616 -628 -597
rect -404 -427 -370 -408
rect -404 -495 -370 -493
rect -404 -531 -370 -529
rect -404 -616 -370 -597
rect -146 -427 -112 -408
rect -146 -495 -112 -493
rect -146 -531 -112 -529
rect -146 -616 -112 -597
rect 112 -427 146 -408
rect 112 -495 146 -493
rect 112 -531 146 -529
rect 112 -616 146 -597
rect 370 -427 404 -408
rect 370 -495 404 -493
rect 370 -531 404 -529
rect 370 -616 404 -597
rect 628 -427 662 -408
rect 628 -495 662 -493
rect 628 -531 662 -529
rect 628 -616 662 -597
rect 886 -427 920 -408
rect 886 -495 920 -493
rect 886 -531 920 -529
rect 886 -616 920 -597
rect -874 -693 -827 -659
rect -791 -693 -757 -659
rect -721 -693 -674 -659
rect -616 -693 -569 -659
rect -533 -693 -499 -659
rect -463 -693 -416 -659
rect -358 -693 -311 -659
rect -275 -693 -241 -659
rect -205 -693 -158 -659
rect -100 -693 -53 -659
rect -17 -693 17 -659
rect 53 -693 100 -659
rect 158 -693 205 -659
rect 241 -693 275 -659
rect 311 -693 358 -659
rect 416 -693 463 -659
rect 499 -693 533 -659
rect 569 -693 616 -659
rect 674 -693 721 -659
rect 757 -693 791 -659
rect 827 -693 874 -659
<< viali >>
rect -920 634 -886 636
rect -920 602 -886 634
rect -920 532 -886 564
rect -920 530 -886 532
rect -662 634 -628 636
rect -662 602 -628 634
rect -662 532 -628 564
rect -662 530 -628 532
rect -404 634 -370 636
rect -404 602 -370 634
rect -404 532 -370 564
rect -404 530 -370 532
rect -146 634 -112 636
rect -146 602 -112 634
rect -146 532 -112 564
rect -146 530 -112 532
rect 112 634 146 636
rect 112 602 146 634
rect 112 532 146 564
rect 112 530 146 532
rect 370 634 404 636
rect 370 602 404 634
rect 370 532 404 564
rect 370 530 404 532
rect 628 634 662 636
rect 628 602 662 634
rect 628 532 662 564
rect 628 530 662 532
rect 886 634 920 636
rect 886 602 920 634
rect 886 532 920 564
rect 886 530 920 532
rect -827 402 -825 436
rect -825 402 -793 436
rect -755 402 -723 436
rect -723 402 -721 436
rect -569 402 -567 436
rect -567 402 -535 436
rect -497 402 -465 436
rect -465 402 -463 436
rect -311 402 -309 436
rect -309 402 -277 436
rect -239 402 -207 436
rect -207 402 -205 436
rect -53 402 -51 436
rect -51 402 -19 436
rect 19 402 51 436
rect 51 402 53 436
rect 205 402 207 436
rect 207 402 239 436
rect 277 402 309 436
rect 309 402 311 436
rect 463 402 465 436
rect 465 402 497 436
rect 535 402 567 436
rect 567 402 569 436
rect 721 402 723 436
rect 723 402 755 436
rect 793 402 825 436
rect 825 402 827 436
rect -920 269 -886 271
rect -920 237 -886 269
rect -920 167 -886 199
rect -920 165 -886 167
rect -662 269 -628 271
rect -662 237 -628 269
rect -662 167 -628 199
rect -662 165 -628 167
rect -404 269 -370 271
rect -404 237 -370 269
rect -404 167 -370 199
rect -404 165 -370 167
rect -146 269 -112 271
rect -146 237 -112 269
rect -146 167 -112 199
rect -146 165 -112 167
rect 112 269 146 271
rect 112 237 146 269
rect 112 167 146 199
rect 112 165 146 167
rect 370 269 404 271
rect 370 237 404 269
rect 370 167 404 199
rect 370 165 404 167
rect 628 269 662 271
rect 628 237 662 269
rect 628 167 662 199
rect 628 165 662 167
rect 886 269 920 271
rect 886 237 920 269
rect 886 167 920 199
rect 886 165 920 167
rect -827 37 -825 71
rect -825 37 -793 71
rect -755 37 -723 71
rect -723 37 -721 71
rect -569 37 -567 71
rect -567 37 -535 71
rect -497 37 -465 71
rect -465 37 -463 71
rect -311 37 -309 71
rect -309 37 -277 71
rect -239 37 -207 71
rect -207 37 -205 71
rect -53 37 -51 71
rect -51 37 -19 71
rect 19 37 51 71
rect 51 37 53 71
rect 205 37 207 71
rect 207 37 239 71
rect 277 37 309 71
rect 309 37 311 71
rect 463 37 465 71
rect 465 37 497 71
rect 535 37 567 71
rect 567 37 569 71
rect 721 37 723 71
rect 723 37 755 71
rect 793 37 825 71
rect 825 37 827 71
rect -920 -96 -886 -94
rect -920 -128 -886 -96
rect -920 -198 -886 -166
rect -920 -200 -886 -198
rect -662 -96 -628 -94
rect -662 -128 -628 -96
rect -662 -198 -628 -166
rect -662 -200 -628 -198
rect -404 -96 -370 -94
rect -404 -128 -370 -96
rect -404 -198 -370 -166
rect -404 -200 -370 -198
rect -146 -96 -112 -94
rect -146 -128 -112 -96
rect -146 -198 -112 -166
rect -146 -200 -112 -198
rect 112 -96 146 -94
rect 112 -128 146 -96
rect 112 -198 146 -166
rect 112 -200 146 -198
rect 370 -96 404 -94
rect 370 -128 404 -96
rect 370 -198 404 -166
rect 370 -200 404 -198
rect 628 -96 662 -94
rect 628 -128 662 -96
rect 628 -198 662 -166
rect 628 -200 662 -198
rect 886 -96 920 -94
rect 886 -128 920 -96
rect 886 -198 920 -166
rect 886 -200 920 -198
rect -827 -328 -825 -294
rect -825 -328 -793 -294
rect -755 -328 -723 -294
rect -723 -328 -721 -294
rect -569 -328 -567 -294
rect -567 -328 -535 -294
rect -497 -328 -465 -294
rect -465 -328 -463 -294
rect -311 -328 -309 -294
rect -309 -328 -277 -294
rect -239 -328 -207 -294
rect -207 -328 -205 -294
rect -53 -328 -51 -294
rect -51 -328 -19 -294
rect 19 -328 51 -294
rect 51 -328 53 -294
rect 205 -328 207 -294
rect 207 -328 239 -294
rect 277 -328 309 -294
rect 309 -328 311 -294
rect 463 -328 465 -294
rect 465 -328 497 -294
rect 535 -328 567 -294
rect 567 -328 569 -294
rect 721 -328 723 -294
rect 723 -328 755 -294
rect 793 -328 825 -294
rect 825 -328 827 -294
rect -920 -461 -886 -459
rect -920 -493 -886 -461
rect -920 -563 -886 -531
rect -920 -565 -886 -563
rect -662 -461 -628 -459
rect -662 -493 -628 -461
rect -662 -563 -628 -531
rect -662 -565 -628 -563
rect -404 -461 -370 -459
rect -404 -493 -370 -461
rect -404 -563 -370 -531
rect -404 -565 -370 -563
rect -146 -461 -112 -459
rect -146 -493 -112 -461
rect -146 -563 -112 -531
rect -146 -565 -112 -563
rect 112 -461 146 -459
rect 112 -493 146 -461
rect 112 -563 146 -531
rect 112 -565 146 -563
rect 370 -461 404 -459
rect 370 -493 404 -461
rect 370 -563 404 -531
rect 370 -565 404 -563
rect 628 -461 662 -459
rect 628 -493 662 -461
rect 628 -563 662 -531
rect 628 -565 662 -563
rect 886 -461 920 -459
rect 886 -493 920 -461
rect 886 -563 920 -531
rect 886 -565 920 -563
rect -827 -693 -825 -659
rect -825 -693 -793 -659
rect -755 -693 -723 -659
rect -723 -693 -721 -659
rect -569 -693 -567 -659
rect -567 -693 -535 -659
rect -497 -693 -465 -659
rect -465 -693 -463 -659
rect -311 -693 -309 -659
rect -309 -693 -277 -659
rect -239 -693 -207 -659
rect -207 -693 -205 -659
rect -53 -693 -51 -659
rect -51 -693 -19 -659
rect 19 -693 51 -659
rect 51 -693 53 -659
rect 205 -693 207 -659
rect 207 -693 239 -659
rect 277 -693 309 -659
rect 309 -693 311 -659
rect 463 -693 465 -659
rect 465 -693 497 -659
rect 535 -693 567 -659
rect 567 -693 569 -659
rect 721 -693 723 -659
rect 723 -693 755 -659
rect 793 -693 825 -659
rect 825 -693 827 -659
<< metal1 >>
rect -926 636 -880 683
rect -926 602 -920 636
rect -886 602 -880 636
rect -926 564 -880 602
rect -926 530 -920 564
rect -886 530 -880 564
rect -926 483 -880 530
rect -668 636 -622 683
rect -668 602 -662 636
rect -628 602 -622 636
rect -668 564 -622 602
rect -668 530 -662 564
rect -628 530 -622 564
rect -668 483 -622 530
rect -410 636 -364 683
rect -410 602 -404 636
rect -370 602 -364 636
rect -410 564 -364 602
rect -410 530 -404 564
rect -370 530 -364 564
rect -410 483 -364 530
rect -152 636 -106 683
rect -152 602 -146 636
rect -112 602 -106 636
rect -152 564 -106 602
rect -152 530 -146 564
rect -112 530 -106 564
rect -152 483 -106 530
rect 106 636 152 683
rect 106 602 112 636
rect 146 602 152 636
rect 106 564 152 602
rect 106 530 112 564
rect 146 530 152 564
rect 106 483 152 530
rect 364 636 410 683
rect 364 602 370 636
rect 404 602 410 636
rect 364 564 410 602
rect 364 530 370 564
rect 404 530 410 564
rect 364 483 410 530
rect 622 636 668 683
rect 622 602 628 636
rect 662 602 668 636
rect 622 564 668 602
rect 622 530 628 564
rect 662 530 668 564
rect 622 483 668 530
rect 880 636 926 683
rect 880 602 886 636
rect 920 602 926 636
rect 880 564 926 602
rect 880 530 886 564
rect 920 530 926 564
rect 880 483 926 530
rect -870 436 -678 442
rect -870 402 -827 436
rect -793 402 -755 436
rect -721 402 -678 436
rect -870 396 -678 402
rect -612 436 -420 442
rect -612 402 -569 436
rect -535 402 -497 436
rect -463 402 -420 436
rect -612 396 -420 402
rect -354 436 -162 442
rect -354 402 -311 436
rect -277 402 -239 436
rect -205 402 -162 436
rect -354 396 -162 402
rect -96 436 96 442
rect -96 402 -53 436
rect -19 402 19 436
rect 53 402 96 436
rect -96 396 96 402
rect 162 436 354 442
rect 162 402 205 436
rect 239 402 277 436
rect 311 402 354 436
rect 162 396 354 402
rect 420 436 612 442
rect 420 402 463 436
rect 497 402 535 436
rect 569 402 612 436
rect 420 396 612 402
rect 678 436 870 442
rect 678 402 721 436
rect 755 402 793 436
rect 827 402 870 436
rect 678 396 870 402
rect -926 271 -880 318
rect -926 237 -920 271
rect -886 237 -880 271
rect -926 199 -880 237
rect -926 165 -920 199
rect -886 165 -880 199
rect -926 118 -880 165
rect -668 271 -622 318
rect -668 237 -662 271
rect -628 237 -622 271
rect -668 199 -622 237
rect -668 165 -662 199
rect -628 165 -622 199
rect -668 118 -622 165
rect -410 271 -364 318
rect -410 237 -404 271
rect -370 237 -364 271
rect -410 199 -364 237
rect -410 165 -404 199
rect -370 165 -364 199
rect -410 118 -364 165
rect -152 271 -106 318
rect -152 237 -146 271
rect -112 237 -106 271
rect -152 199 -106 237
rect -152 165 -146 199
rect -112 165 -106 199
rect -152 118 -106 165
rect 106 271 152 318
rect 106 237 112 271
rect 146 237 152 271
rect 106 199 152 237
rect 106 165 112 199
rect 146 165 152 199
rect 106 118 152 165
rect 364 271 410 318
rect 364 237 370 271
rect 404 237 410 271
rect 364 199 410 237
rect 364 165 370 199
rect 404 165 410 199
rect 364 118 410 165
rect 622 271 668 318
rect 622 237 628 271
rect 662 237 668 271
rect 622 199 668 237
rect 622 165 628 199
rect 662 165 668 199
rect 622 118 668 165
rect 880 271 926 318
rect 880 237 886 271
rect 920 237 926 271
rect 880 199 926 237
rect 880 165 886 199
rect 920 165 926 199
rect 880 118 926 165
rect -870 71 -678 77
rect -870 37 -827 71
rect -793 37 -755 71
rect -721 37 -678 71
rect -870 31 -678 37
rect -612 71 -420 77
rect -612 37 -569 71
rect -535 37 -497 71
rect -463 37 -420 71
rect -612 31 -420 37
rect -354 71 -162 77
rect -354 37 -311 71
rect -277 37 -239 71
rect -205 37 -162 71
rect -354 31 -162 37
rect -96 71 96 77
rect -96 37 -53 71
rect -19 37 19 71
rect 53 37 96 71
rect -96 31 96 37
rect 162 71 354 77
rect 162 37 205 71
rect 239 37 277 71
rect 311 37 354 71
rect 162 31 354 37
rect 420 71 612 77
rect 420 37 463 71
rect 497 37 535 71
rect 569 37 612 71
rect 420 31 612 37
rect 678 71 870 77
rect 678 37 721 71
rect 755 37 793 71
rect 827 37 870 71
rect 678 31 870 37
rect -926 -94 -880 -47
rect -926 -128 -920 -94
rect -886 -128 -880 -94
rect -926 -166 -880 -128
rect -926 -200 -920 -166
rect -886 -200 -880 -166
rect -926 -247 -880 -200
rect -668 -94 -622 -47
rect -668 -128 -662 -94
rect -628 -128 -622 -94
rect -668 -166 -622 -128
rect -668 -200 -662 -166
rect -628 -200 -622 -166
rect -668 -247 -622 -200
rect -410 -94 -364 -47
rect -410 -128 -404 -94
rect -370 -128 -364 -94
rect -410 -166 -364 -128
rect -410 -200 -404 -166
rect -370 -200 -364 -166
rect -410 -247 -364 -200
rect -152 -94 -106 -47
rect -152 -128 -146 -94
rect -112 -128 -106 -94
rect -152 -166 -106 -128
rect -152 -200 -146 -166
rect -112 -200 -106 -166
rect -152 -247 -106 -200
rect 106 -94 152 -47
rect 106 -128 112 -94
rect 146 -128 152 -94
rect 106 -166 152 -128
rect 106 -200 112 -166
rect 146 -200 152 -166
rect 106 -247 152 -200
rect 364 -94 410 -47
rect 364 -128 370 -94
rect 404 -128 410 -94
rect 364 -166 410 -128
rect 364 -200 370 -166
rect 404 -200 410 -166
rect 364 -247 410 -200
rect 622 -94 668 -47
rect 622 -128 628 -94
rect 662 -128 668 -94
rect 622 -166 668 -128
rect 622 -200 628 -166
rect 662 -200 668 -166
rect 622 -247 668 -200
rect 880 -94 926 -47
rect 880 -128 886 -94
rect 920 -128 926 -94
rect 880 -166 926 -128
rect 880 -200 886 -166
rect 920 -200 926 -166
rect 880 -247 926 -200
rect -870 -294 -678 -288
rect -870 -328 -827 -294
rect -793 -328 -755 -294
rect -721 -328 -678 -294
rect -870 -334 -678 -328
rect -612 -294 -420 -288
rect -612 -328 -569 -294
rect -535 -328 -497 -294
rect -463 -328 -420 -294
rect -612 -334 -420 -328
rect -354 -294 -162 -288
rect -354 -328 -311 -294
rect -277 -328 -239 -294
rect -205 -328 -162 -294
rect -354 -334 -162 -328
rect -96 -294 96 -288
rect -96 -328 -53 -294
rect -19 -328 19 -294
rect 53 -328 96 -294
rect -96 -334 96 -328
rect 162 -294 354 -288
rect 162 -328 205 -294
rect 239 -328 277 -294
rect 311 -328 354 -294
rect 162 -334 354 -328
rect 420 -294 612 -288
rect 420 -328 463 -294
rect 497 -328 535 -294
rect 569 -328 612 -294
rect 420 -334 612 -328
rect 678 -294 870 -288
rect 678 -328 721 -294
rect 755 -328 793 -294
rect 827 -328 870 -294
rect 678 -334 870 -328
rect -926 -459 -880 -412
rect -926 -493 -920 -459
rect -886 -493 -880 -459
rect -926 -531 -880 -493
rect -926 -565 -920 -531
rect -886 -565 -880 -531
rect -926 -612 -880 -565
rect -668 -459 -622 -412
rect -668 -493 -662 -459
rect -628 -493 -622 -459
rect -668 -531 -622 -493
rect -668 -565 -662 -531
rect -628 -565 -622 -531
rect -668 -612 -622 -565
rect -410 -459 -364 -412
rect -410 -493 -404 -459
rect -370 -493 -364 -459
rect -410 -531 -364 -493
rect -410 -565 -404 -531
rect -370 -565 -364 -531
rect -410 -612 -364 -565
rect -152 -459 -106 -412
rect -152 -493 -146 -459
rect -112 -493 -106 -459
rect -152 -531 -106 -493
rect -152 -565 -146 -531
rect -112 -565 -106 -531
rect -152 -612 -106 -565
rect 106 -459 152 -412
rect 106 -493 112 -459
rect 146 -493 152 -459
rect 106 -531 152 -493
rect 106 -565 112 -531
rect 146 -565 152 -531
rect 106 -612 152 -565
rect 364 -459 410 -412
rect 364 -493 370 -459
rect 404 -493 410 -459
rect 364 -531 410 -493
rect 364 -565 370 -531
rect 404 -565 410 -531
rect 364 -612 410 -565
rect 622 -459 668 -412
rect 622 -493 628 -459
rect 662 -493 668 -459
rect 622 -531 668 -493
rect 622 -565 628 -531
rect 662 -565 668 -531
rect 622 -612 668 -565
rect 880 -459 926 -412
rect 880 -493 886 -459
rect 920 -493 926 -459
rect 880 -531 926 -493
rect 880 -565 886 -531
rect 920 -565 926 -531
rect 880 -612 926 -565
rect -870 -659 -678 -653
rect -870 -693 -827 -659
rect -793 -693 -755 -659
rect -721 -693 -678 -659
rect -870 -699 -678 -693
rect -612 -659 -420 -653
rect -612 -693 -569 -659
rect -535 -693 -497 -659
rect -463 -693 -420 -659
rect -612 -699 -420 -693
rect -354 -659 -162 -653
rect -354 -693 -311 -659
rect -277 -693 -239 -659
rect -205 -693 -162 -659
rect -354 -699 -162 -693
rect -96 -659 96 -653
rect -96 -693 -53 -659
rect -19 -693 19 -659
rect 53 -693 96 -659
rect -96 -699 96 -693
rect 162 -659 354 -653
rect 162 -693 205 -659
rect 239 -693 277 -659
rect 311 -693 354 -659
rect 162 -699 354 -693
rect 420 -659 612 -653
rect 420 -693 463 -659
rect 497 -693 535 -659
rect 569 -693 612 -659
rect 420 -699 612 -693
rect 678 -659 870 -653
rect 678 -693 721 -659
rect 755 -693 793 -659
rect 827 -693 870 -659
rect 678 -699 870 -693
<< end >>
