magic
tech sky130A
timestamp 1662947835
<< metal1 >>
rect -12000 7500 110000 12000
rect -12000 4500 500 7500
rect 99500 4500 110000 7500
rect -12000 -1500 110000 4500
rect -12000 -4500 500 -1500
rect 99500 -4500 110000 -1500
rect -12000 -9000 110000 -4500
rect -12000 -39000 0 -9000
rect 100000 -39000 110000 -9000
rect -12000 -45500 110000 -39000
rect -12000 -48500 500 -45500
rect 99500 -48500 110000 -45500
rect -12000 -54500 110000 -48500
rect -12000 -57500 500 -54500
rect 99500 -57500 110000 -54500
rect -12000 -64000 110000 -57500
<< via1 >>
rect 500 4500 99500 7500
rect 500 -4500 99500 -1500
rect 500 -48500 99500 -45500
rect 500 -57500 99500 -54500
<< metal2 >>
rect 0 7500 100000 8000
rect 0 4500 500 7500
rect 99500 4500 100000 7500
rect 0 4000 100000 4500
rect -1000 1900 101000 2000
rect -1000 1100 -900 1900
rect -100 1100 100100 1900
rect 100900 1100 101000 1900
rect -1000 1000 101000 1100
rect 0 -1500 100000 -1000
rect 0 -4500 500 -1500
rect 99500 -4500 100000 -1500
rect 0 -5000 100000 -4500
rect 0 -45500 100000 -45000
rect 0 -48500 500 -45500
rect 99500 -48500 100000 -45500
rect 0 -49000 100000 -48500
rect -1000 -51100 101000 -51000
rect -1000 -51900 -900 -51100
rect -100 -51900 100100 -51100
rect 100900 -51900 101000 -51100
rect -1000 -52000 101000 -51900
rect 0 -54500 100000 -54000
rect 0 -57500 500 -54500
rect 99500 -57500 100000 -54500
rect 0 -58000 100000 -57500
<< via2 >>
rect -900 1100 -100 1900
rect 100100 1100 100900 1900
rect -900 -51900 -100 -51100
rect 100100 -51900 100900 -51100
<< metal3 >>
rect -1000 1900 0 2000
rect -1000 1100 -900 1900
rect -100 1100 0 1900
rect -1000 1000 0 1100
rect 100000 1900 101000 2000
rect 100000 1100 100100 1900
rect 100900 1100 101000 1900
rect 100000 1000 101000 1100
rect -1000 -51100 0 -51000
rect -1000 -51900 -900 -51100
rect -100 -51900 0 -51100
rect -1000 -52000 0 -51900
rect 100000 -51100 101000 -51000
rect 100000 -51900 100100 -51100
rect 100900 -51900 101000 -51100
rect 100000 -52000 101000 -51900
<< labels >>
flabel metal3 -1000 1000 -900 2000 0 FreeSans 20000 0 0 0 INA
flabel metal3 -1000 -52000 -900 -51000 0 FreeSans 20000 0 0 0 INB
flabel metal3 100900 1000 101000 2000 0 FreeSans 20000 0 0 0 OUTA
flabel metal3 100900 -52000 101000 -51000 0 FreeSans 20000 0 0 0 OUTB
flabel metal1 -12000 -64000 110000 -57500 0 FreeSans 20000 0 0 0 GND
<< end >>
