magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -297 2102 297 2188
rect -297 -2102 -211 2102
rect 211 -2102 297 2102
rect -297 -2188 297 -2102
<< psubdiff >>
rect -271 2128 -153 2162
rect -119 2128 -85 2162
rect -51 2128 -17 2162
rect 17 2128 51 2162
rect 85 2128 119 2162
rect 153 2128 271 2162
rect -271 2057 -237 2128
rect 237 2057 271 2128
rect -271 1989 -237 2023
rect -271 1921 -237 1955
rect -271 1853 -237 1887
rect -271 1785 -237 1819
rect -271 1717 -237 1751
rect -271 1649 -237 1683
rect -271 1581 -237 1615
rect -271 1513 -237 1547
rect -271 1445 -237 1479
rect -271 1377 -237 1411
rect -271 1309 -237 1343
rect -271 1241 -237 1275
rect -271 1173 -237 1207
rect -271 1105 -237 1139
rect -271 1037 -237 1071
rect -271 969 -237 1003
rect -271 901 -237 935
rect -271 833 -237 867
rect -271 765 -237 799
rect -271 697 -237 731
rect -271 629 -237 663
rect -271 561 -237 595
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect -271 -595 -237 -561
rect -271 -663 -237 -629
rect -271 -731 -237 -697
rect -271 -799 -237 -765
rect -271 -867 -237 -833
rect -271 -935 -237 -901
rect -271 -1003 -237 -969
rect -271 -1071 -237 -1037
rect -271 -1139 -237 -1105
rect -271 -1207 -237 -1173
rect -271 -1275 -237 -1241
rect -271 -1343 -237 -1309
rect -271 -1411 -237 -1377
rect -271 -1479 -237 -1445
rect -271 -1547 -237 -1513
rect -271 -1615 -237 -1581
rect -271 -1683 -237 -1649
rect -271 -1751 -237 -1717
rect -271 -1819 -237 -1785
rect -271 -1887 -237 -1853
rect -271 -1955 -237 -1921
rect -271 -2023 -237 -1989
rect 237 1989 271 2023
rect 237 1921 271 1955
rect 237 1853 271 1887
rect 237 1785 271 1819
rect 237 1717 271 1751
rect 237 1649 271 1683
rect 237 1581 271 1615
rect 237 1513 271 1547
rect 237 1445 271 1479
rect 237 1377 271 1411
rect 237 1309 271 1343
rect 237 1241 271 1275
rect 237 1173 271 1207
rect 237 1105 271 1139
rect 237 1037 271 1071
rect 237 969 271 1003
rect 237 901 271 935
rect 237 833 271 867
rect 237 765 271 799
rect 237 697 271 731
rect 237 629 271 663
rect 237 561 271 595
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect 237 -595 271 -561
rect 237 -663 271 -629
rect 237 -731 271 -697
rect 237 -799 271 -765
rect 237 -867 271 -833
rect 237 -935 271 -901
rect 237 -1003 271 -969
rect 237 -1071 271 -1037
rect 237 -1139 271 -1105
rect 237 -1207 271 -1173
rect 237 -1275 271 -1241
rect 237 -1343 271 -1309
rect 237 -1411 271 -1377
rect 237 -1479 271 -1445
rect 237 -1547 271 -1513
rect 237 -1615 271 -1581
rect 237 -1683 271 -1649
rect 237 -1751 271 -1717
rect 237 -1819 271 -1785
rect 237 -1887 271 -1853
rect 237 -1955 271 -1921
rect 237 -2023 271 -1989
rect -271 -2128 -237 -2057
rect 237 -2128 271 -2057
rect -271 -2162 -153 -2128
rect -119 -2162 -85 -2128
rect -51 -2162 -17 -2128
rect 17 -2162 51 -2128
rect 85 -2162 119 -2128
rect 153 -2162 271 -2128
<< psubdiffcont >>
rect -153 2128 -119 2162
rect -85 2128 -51 2162
rect -17 2128 17 2162
rect 51 2128 85 2162
rect 119 2128 153 2162
rect -271 2023 -237 2057
rect -271 1955 -237 1989
rect -271 1887 -237 1921
rect -271 1819 -237 1853
rect -271 1751 -237 1785
rect -271 1683 -237 1717
rect -271 1615 -237 1649
rect -271 1547 -237 1581
rect -271 1479 -237 1513
rect -271 1411 -237 1445
rect -271 1343 -237 1377
rect -271 1275 -237 1309
rect -271 1207 -237 1241
rect -271 1139 -237 1173
rect -271 1071 -237 1105
rect -271 1003 -237 1037
rect -271 935 -237 969
rect -271 867 -237 901
rect -271 799 -237 833
rect -271 731 -237 765
rect -271 663 -237 697
rect -271 595 -237 629
rect -271 527 -237 561
rect -271 459 -237 493
rect -271 391 -237 425
rect -271 323 -237 357
rect -271 255 -237 289
rect -271 187 -237 221
rect -271 119 -237 153
rect -271 51 -237 85
rect -271 -17 -237 17
rect -271 -85 -237 -51
rect -271 -153 -237 -119
rect -271 -221 -237 -187
rect -271 -289 -237 -255
rect -271 -357 -237 -323
rect -271 -425 -237 -391
rect -271 -493 -237 -459
rect -271 -561 -237 -527
rect -271 -629 -237 -595
rect -271 -697 -237 -663
rect -271 -765 -237 -731
rect -271 -833 -237 -799
rect -271 -901 -237 -867
rect -271 -969 -237 -935
rect -271 -1037 -237 -1003
rect -271 -1105 -237 -1071
rect -271 -1173 -237 -1139
rect -271 -1241 -237 -1207
rect -271 -1309 -237 -1275
rect -271 -1377 -237 -1343
rect -271 -1445 -237 -1411
rect -271 -1513 -237 -1479
rect -271 -1581 -237 -1547
rect -271 -1649 -237 -1615
rect -271 -1717 -237 -1683
rect -271 -1785 -237 -1751
rect -271 -1853 -237 -1819
rect -271 -1921 -237 -1887
rect -271 -1989 -237 -1955
rect -271 -2057 -237 -2023
rect 237 2023 271 2057
rect 237 1955 271 1989
rect 237 1887 271 1921
rect 237 1819 271 1853
rect 237 1751 271 1785
rect 237 1683 271 1717
rect 237 1615 271 1649
rect 237 1547 271 1581
rect 237 1479 271 1513
rect 237 1411 271 1445
rect 237 1343 271 1377
rect 237 1275 271 1309
rect 237 1207 271 1241
rect 237 1139 271 1173
rect 237 1071 271 1105
rect 237 1003 271 1037
rect 237 935 271 969
rect 237 867 271 901
rect 237 799 271 833
rect 237 731 271 765
rect 237 663 271 697
rect 237 595 271 629
rect 237 527 271 561
rect 237 459 271 493
rect 237 391 271 425
rect 237 323 271 357
rect 237 255 271 289
rect 237 187 271 221
rect 237 119 271 153
rect 237 51 271 85
rect 237 -17 271 17
rect 237 -85 271 -51
rect 237 -153 271 -119
rect 237 -221 271 -187
rect 237 -289 271 -255
rect 237 -357 271 -323
rect 237 -425 271 -391
rect 237 -493 271 -459
rect 237 -561 271 -527
rect 237 -629 271 -595
rect 237 -697 271 -663
rect 237 -765 271 -731
rect 237 -833 271 -799
rect 237 -901 271 -867
rect 237 -969 271 -935
rect 237 -1037 271 -1003
rect 237 -1105 271 -1071
rect 237 -1173 271 -1139
rect 237 -1241 271 -1207
rect 237 -1309 271 -1275
rect 237 -1377 271 -1343
rect 237 -1445 271 -1411
rect 237 -1513 271 -1479
rect 237 -1581 271 -1547
rect 237 -1649 271 -1615
rect 237 -1717 271 -1683
rect 237 -1785 271 -1751
rect 237 -1853 271 -1819
rect 237 -1921 271 -1887
rect 237 -1989 271 -1955
rect 237 -2057 271 -2023
rect -153 -2162 -119 -2128
rect -85 -2162 -51 -2128
rect -17 -2162 17 -2128
rect 51 -2162 85 -2128
rect 119 -2162 153 -2128
<< xpolycontact >>
rect -141 1600 141 2032
rect -141 -2032 141 -1600
<< ppolyres >>
rect -141 -1600 141 1600
<< locali >>
rect -271 2128 -153 2162
rect -119 2128 -85 2162
rect -51 2128 -17 2162
rect 17 2128 51 2162
rect 85 2128 119 2162
rect 153 2128 271 2162
rect -271 2057 -237 2128
rect 237 2057 271 2128
rect -271 1989 -237 2023
rect -271 1921 -237 1955
rect -271 1853 -237 1887
rect -271 1785 -237 1819
rect -271 1717 -237 1751
rect -271 1649 -237 1683
rect -271 1581 -237 1615
rect 237 1989 271 2023
rect 237 1921 271 1955
rect 237 1853 271 1887
rect 237 1785 271 1819
rect 237 1717 271 1751
rect 237 1649 271 1683
rect -271 1513 -237 1547
rect -271 1445 -237 1479
rect -271 1377 -237 1411
rect -271 1309 -237 1343
rect -271 1241 -237 1275
rect -271 1173 -237 1207
rect -271 1105 -237 1139
rect -271 1037 -237 1071
rect -271 969 -237 1003
rect -271 901 -237 935
rect -271 833 -237 867
rect -271 765 -237 799
rect -271 697 -237 731
rect -271 629 -237 663
rect -271 561 -237 595
rect -271 493 -237 527
rect -271 425 -237 459
rect -271 357 -237 391
rect -271 289 -237 323
rect -271 221 -237 255
rect -271 153 -237 187
rect -271 85 -237 119
rect -271 17 -237 51
rect -271 -51 -237 -17
rect -271 -119 -237 -85
rect -271 -187 -237 -153
rect -271 -255 -237 -221
rect -271 -323 -237 -289
rect -271 -391 -237 -357
rect -271 -459 -237 -425
rect -271 -527 -237 -493
rect -271 -595 -237 -561
rect -271 -663 -237 -629
rect -271 -731 -237 -697
rect -271 -799 -237 -765
rect -271 -867 -237 -833
rect -271 -935 -237 -901
rect -271 -1003 -237 -969
rect -271 -1071 -237 -1037
rect -271 -1139 -237 -1105
rect -271 -1207 -237 -1173
rect -271 -1275 -237 -1241
rect -271 -1343 -237 -1309
rect -271 -1411 -237 -1377
rect -271 -1479 -237 -1445
rect -271 -1547 -237 -1513
rect -271 -1615 -237 -1581
rect 237 1581 271 1615
rect 237 1513 271 1547
rect 237 1445 271 1479
rect 237 1377 271 1411
rect 237 1309 271 1343
rect 237 1241 271 1275
rect 237 1173 271 1207
rect 237 1105 271 1139
rect 237 1037 271 1071
rect 237 969 271 1003
rect 237 901 271 935
rect 237 833 271 867
rect 237 765 271 799
rect 237 697 271 731
rect 237 629 271 663
rect 237 561 271 595
rect 237 493 271 527
rect 237 425 271 459
rect 237 357 271 391
rect 237 289 271 323
rect 237 221 271 255
rect 237 153 271 187
rect 237 85 271 119
rect 237 17 271 51
rect 237 -51 271 -17
rect 237 -119 271 -85
rect 237 -187 271 -153
rect 237 -255 271 -221
rect 237 -323 271 -289
rect 237 -391 271 -357
rect 237 -459 271 -425
rect 237 -527 271 -493
rect 237 -595 271 -561
rect 237 -663 271 -629
rect 237 -731 271 -697
rect 237 -799 271 -765
rect 237 -867 271 -833
rect 237 -935 271 -901
rect 237 -1003 271 -969
rect 237 -1071 271 -1037
rect 237 -1139 271 -1105
rect 237 -1207 271 -1173
rect 237 -1275 271 -1241
rect 237 -1343 271 -1309
rect 237 -1411 271 -1377
rect 237 -1479 271 -1445
rect 237 -1547 271 -1513
rect -271 -1683 -237 -1649
rect -271 -1751 -237 -1717
rect -271 -1819 -237 -1785
rect -271 -1887 -237 -1853
rect -271 -1955 -237 -1921
rect -271 -2023 -237 -1989
rect 237 -1615 271 -1581
rect 237 -1683 271 -1649
rect 237 -1751 271 -1717
rect 237 -1819 271 -1785
rect 237 -1887 271 -1853
rect 237 -1955 271 -1921
rect 237 -2023 271 -1989
rect -271 -2128 -237 -2057
rect 237 -2128 271 -2057
rect -271 -2162 -153 -2128
rect -119 -2162 -85 -2128
rect -51 -2162 -17 -2128
rect 17 -2162 51 -2128
rect 85 -2162 119 -2128
rect 153 -2162 271 -2128
<< viali >>
rect -125 1618 125 2012
rect -125 -2013 125 -1619
<< metal1 >>
rect -131 2012 131 2026
rect -131 1618 -125 2012
rect 125 1618 131 2012
rect -131 1605 131 1618
rect -131 -1619 131 -1605
rect -131 -2013 -125 -1619
rect 125 -2013 131 -1619
rect -131 -2026 131 -2013
<< properties >>
string FIXED_BBOX -254 -2145 254 2145
<< end >>
