magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -125 -138 -67 -132
rect 67 -138 125 -132
rect -125 -172 -113 -138
rect 67 -172 79 -138
rect -125 -178 -67 -172
rect 67 -178 125 -172
<< pwell >>
rect -301 -300 301 300
<< nmoslvt >>
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
<< ndiff >>
rect -173 85 -111 100
rect -173 51 -161 85
rect -127 51 -111 85
rect -173 17 -111 51
rect -173 -17 -161 17
rect -127 -17 -111 17
rect -173 -51 -111 -17
rect -173 -85 -161 -51
rect -127 -85 -111 -51
rect -173 -100 -111 -85
rect -81 85 -15 100
rect -81 51 -65 85
rect -31 51 -15 85
rect -81 17 -15 51
rect -81 -17 -65 17
rect -31 -17 -15 17
rect -81 -51 -15 -17
rect -81 -85 -65 -51
rect -31 -85 -15 -51
rect -81 -100 -15 -85
rect 15 85 81 100
rect 15 51 31 85
rect 65 51 81 85
rect 15 17 81 51
rect 15 -17 31 17
rect 65 -17 81 17
rect 15 -51 81 -17
rect 15 -85 31 -51
rect 65 -85 81 -51
rect 15 -100 81 -85
rect 111 85 173 100
rect 111 51 127 85
rect 161 51 173 85
rect 111 17 173 51
rect 111 -17 127 17
rect 161 -17 173 17
rect 111 -51 173 -17
rect 111 -85 127 -51
rect 161 -85 173 -51
rect 111 -100 173 -85
<< ndiffc >>
rect -161 51 -127 85
rect -161 -17 -127 17
rect -161 -85 -127 -51
rect -65 51 -31 85
rect -65 -17 -31 17
rect -65 -85 -31 -51
rect 31 51 65 85
rect 31 -17 65 17
rect 31 -85 65 -51
rect 127 51 161 85
rect 127 -17 161 17
rect 127 -85 161 -51
<< psubdiff >>
rect -275 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 275 274
rect -275 153 -241 240
rect -275 85 -241 119
rect 241 153 275 240
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect -275 -240 -241 -153
rect 241 -119 275 -85
rect 241 -240 275 -153
rect -275 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 275 -240
<< psubdiffcont >>
rect -153 240 -119 274
rect -85 240 -51 274
rect -17 240 17 274
rect 51 240 85 274
rect 119 240 153 274
rect -275 119 -241 153
rect 241 119 275 153
rect -275 51 -241 85
rect -275 -17 -241 17
rect -275 -85 -241 -51
rect 241 51 275 85
rect 241 -17 275 17
rect 241 -85 275 -51
rect -275 -153 -241 -119
rect 241 -153 275 -119
rect -153 -274 -119 -240
rect -85 -274 -51 -240
rect -17 -274 17 -240
rect 51 -274 85 -240
rect 119 -274 153 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -111 100 -81 126
rect -33 122 33 138
rect -15 100 15 122
rect 81 100 111 126
rect -111 -122 -81 -100
rect -129 -138 -63 -122
rect -15 -126 15 -100
rect 81 -122 111 -100
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect -129 -188 -63 -172
rect 63 -138 129 -122
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 63 -188 129 -172
<< polycont >>
rect -17 138 17 172
rect -113 -172 -79 -138
rect 79 -172 113 -138
<< locali >>
rect -275 240 -153 274
rect -119 240 -85 274
rect -51 240 -17 274
rect 17 240 51 274
rect 85 240 119 274
rect 153 240 275 274
rect -275 153 -241 240
rect -33 138 -17 172
rect 17 138 33 172
rect 241 153 275 240
rect -275 85 -241 119
rect -275 17 -241 51
rect -275 -51 -241 -17
rect -275 -119 -241 -85
rect -161 85 -127 104
rect -161 17 -127 19
rect -161 -19 -127 -17
rect -161 -104 -127 -85
rect -65 85 -31 104
rect -65 17 -31 19
rect -65 -19 -31 -17
rect -65 -104 -31 -85
rect 31 85 65 104
rect 31 17 65 19
rect 31 -19 65 -17
rect 31 -104 65 -85
rect 127 85 161 104
rect 127 17 161 19
rect 127 -19 161 -17
rect 127 -104 161 -85
rect 241 85 275 119
rect 241 17 275 51
rect 241 -51 275 -17
rect 241 -119 275 -85
rect -275 -240 -241 -153
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 241 -240 275 -153
rect -275 -274 -153 -240
rect -119 -274 -85 -240
rect -51 -274 -17 -240
rect 17 -274 51 -240
rect 85 -274 119 -240
rect 153 -274 275 -240
<< viali >>
rect -17 138 17 172
rect -161 51 -127 53
rect -161 19 -127 51
rect -161 -51 -127 -19
rect -161 -53 -127 -51
rect -65 51 -31 53
rect -65 19 -31 51
rect -65 -51 -31 -19
rect -65 -53 -31 -51
rect 31 51 65 53
rect 31 19 65 51
rect 31 -51 65 -19
rect 31 -53 65 -51
rect 127 51 161 53
rect 127 19 161 51
rect 127 -51 161 -19
rect 127 -53 161 -51
rect -113 -172 -79 -138
rect 79 -172 113 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -167 53 -121 100
rect -167 19 -161 53
rect -127 19 -121 53
rect -167 -19 -121 19
rect -167 -53 -161 -19
rect -127 -53 -121 -19
rect -167 -100 -121 -53
rect -71 53 -25 100
rect -71 19 -65 53
rect -31 19 -25 53
rect -71 -19 -25 19
rect -71 -53 -65 -19
rect -31 -53 -25 -19
rect -71 -100 -25 -53
rect 25 53 71 100
rect 25 19 31 53
rect 65 19 71 53
rect 25 -19 71 19
rect 25 -53 31 -19
rect 65 -53 71 -19
rect 25 -100 71 -53
rect 121 53 167 100
rect 121 19 127 53
rect 161 19 167 53
rect 121 -19 167 19
rect 121 -53 127 -19
rect 161 -53 167 -19
rect 121 -100 167 -53
rect -125 -138 -67 -132
rect -125 -172 -113 -138
rect -79 -172 -67 -138
rect -125 -178 -67 -172
rect 67 -138 125 -132
rect 67 -172 79 -138
rect 113 -172 125 -138
rect 67 -178 125 -172
<< properties >>
string FIXED_BBOX -258 -257 258 257
<< end >>
