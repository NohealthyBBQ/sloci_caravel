* NGSPICE file created from user_analog_project_wrapper.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_lvt_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_DJ7QE5 a_15_122# a_n227_n274# a_n125_n100# a_n81_n188#
+ a_63_n100# a_n33_n100#
X0 a_63_n100# a_15_122# a_n33_n100# a_n227_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n188# a_n125_n100# a_n227_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_BX7S53 a_n275_n274# a_n173_n100# a_15_n100# a_n33_122#
+ a_111_n100# a_n81_n100# a_n129_n188# a_63_n188#
X0 a_15_n100# a_n33_122# a_n81_n100# a_n275_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n81_n100# a_n129_n188# a_n173_n100# a_n275_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X2 a_111_n100# a_63_n188# a_15_n100# a_n275_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_B6HS5D a_159_n100# a_111_n188# a_15_122# a_n273_n188#
+ a_255_n100# a_207_122# a_n129_n100# a_n81_n188# a_63_n100# a_n177_122# a_n225_n100#
+ a_n33_n100# a_n419_n274# a_n317_n100#
X0 a_63_n100# a_15_122# a_n33_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n188# a_n129_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_159_n100# a_111_n188# a_63_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_255_n100# a_207_122# a_159_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n225_n100# a_n273_n188# a_n317_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X5 a_n129_n100# a_n177_122# a_n225_n100# a_n419_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_WCTBV5 m4_n551_n300# c2_n451_n200#
X0 c2_n451_n200# m4_n551_n300# sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_WCTZRP c2_n551_n200# m4_n651_n300#
X0 c2_n551_n200# m4_n651_n300# sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=3e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_3ZFDVT c2_n551_n400# m4_n651_n500#
X0 c2_n551_n400# m4_n651_n500# sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=3e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_VCH7EQ c2_n851_n400# m4_n951_n500#
X0 c2_n851_n400# m4_n951_n500# sky130_fd_pr__cap_mim_m3_2 l=4e+06u w=6e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_2_FJFAMD m4_n551_n300# c2_n451_n200#
X0 c2_n451_n200# m4_n551_n300# sky130_fd_pr__cap_mim_m3_2 l=2e+06u w=2e+06u
.ends

.subckt cap_bank ctrll5 ctrll4 ctrll2 ctrll3 ctrll1 IN GND
XXM1 m1_3910_n1320# ctrll1 GND GND sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM2 GND ctrll2 m1_4820_n1420# GND sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM3 ctrll3 GND GND ctrll3 GND m1_4820_n890# sky130_fd_pr__nfet_01v8_lvt_DJ7QE5
XXM4 GND GND GND ctrll4 m1_4820_n460# m1_4820_n460# ctrll4 ctrll4 sky130_fd_pr__nfet_01v8_lvt_BX7S53
XXM5 m1_4700_270# ctrll5 ctrll5 ctrll5 GND ctrll5 GND ctrll5 GND ctrll5 m1_4700_270#
+ m1_4700_270# GND GND sky130_fd_pr__nfet_01v8_lvt_B6HS5D
XXC1 m1_4820_n1420# IN sky130_fd_pr__cap_mim_m3_2_WCTBV5
XXC2 IN m1_4820_n890# sky130_fd_pr__cap_mim_m3_2_WCTZRP
XXC3 IN m1_4820_n460# sky130_fd_pr__cap_mim_m3_2_3ZFDVT
XXC4 IN m1_4700_270# sky130_fd_pr__cap_mim_m3_2_VCH7EQ
XXC6 m1_3910_n1320# IN sky130_fd_pr__cap_mim_m3_2_FJFAMD
.ends

.subckt sky130_fd_pr__res_high_po_2p85_P79JE3 a_n285_n1192# a_n285_760# a_n415_n1322#
X0 a_n285_n1192# a_n285_760# a_n415_n1322# sky130_fd_pr__res_high_po_2p85 l=7.6e+06u
.ends

.subckt sky130_fd_pr__res_high_po_5p73_W59YBA a_n573_1640# a_n573_n2072# a_n703_n2202#
X0 a_n573_n2072# a_n573_1640# a_n703_n2202# sky130_fd_pr__res_high_po_5p73 l=1.64e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_YTLFGX a_543_n100# a_159_n100# a_n609_n100# a_n705_n100#
+ a_255_n100# a_351_n100# a_n417_n100# a_n801_n100# a_n129_n100# a_n513_n100# a_n989_n100#
+ a_63_n100# a_n225_n100# a_n945_n188# a_927_n100# a_n1091_n274# a_n321_n100# a_639_n100#
+ a_735_n100# a_n33_n100# a_n897_n100# a_831_n100# a_447_n100#
X0 a_63_n100# a_n945_n188# a_n33_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_927_n100# a_n945_n188# a_831_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n33_n100# a_n945_n188# a_n129_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_351_n100# a_n945_n188# a_255_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_159_n100# a_n945_n188# a_63_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_255_n100# a_n945_n188# a_159_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X6 a_447_n100# a_n945_n188# a_351_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_543_n100# a_n945_n188# a_447_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_735_n100# a_n945_n188# a_639_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X9 a_831_n100# a_n945_n188# a_735_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_639_n100# a_n945_n188# a_543_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X11 a_n321_n100# a_n945_n188# a_n417_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_n801_n100# a_n945_n188# a_n897_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n705_n100# a_n945_n188# a_n801_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_n513_n100# a_n945_n188# a_n609_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X15 a_n417_n100# a_n945_n188# a_n513_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_n225_n100# a_n945_n188# a_n321_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_n129_n100# a_n945_n188# a_n225_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_n897_n100# a_n945_n188# a_n989_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X19 a_n609_n100# a_n945_n188# a_n705_n100# a_n1091_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_LELFGX a_543_n100# a_n609_n100# a_159_n100# a_1695_n100#
+ a_n2001_122# a_879_122# a_2655_n100# a_n2481_n188# a_n273_122# a_n1953_n100# a_n2097_n188#
+ a_n1569_n100# a_n1521_n188# a_1839_122# a_n2529_n100# a_n1137_n188# a_n705_n100#
+ a_1791_n100# a_n1233_122# a_255_n100# a_975_n188# a_2751_n100# a_2367_n100# a_1407_n100#
+ a_1071_122# a_n1665_n100# a_n2625_n100# a_n2577_122# a_n801_n100# a_351_n100# a_n417_n100#
+ a_2463_n100# a_2079_n100# a_n465_122# a_1503_n100# a_2031_122# a_n1761_n100# a_1119_n100#
+ a_n2721_n100# a_n1377_n100# a_n2337_n100# a_n1425_122# a_n513_n100# a_783_n188#
+ a_n129_n100# a_399_n188# a_2175_n100# a_1263_122# a_1215_n100# a_n1473_n100# a_63_n100#
+ a_1935_n188# a_n2433_n100# a_n1089_n100# a_n2049_n100# a_n2769_122# a_n2909_n100#
+ a_n225_n100# a_2271_n100# a_n657_122# a_n945_n188# a_2223_122# a_927_n100# a_1311_n100#
+ a_n1185_n100# a_n2145_n100# a_495_122# a_n2865_n188# a_n1617_122# a_n3011_n274#
+ a_111_122# a_n321_n100# a_n1905_n188# a_591_n188# a_1455_122# a_639_n100# a_1023_n100#
+ a_207_n188# a_1743_n188# a_n1281_n100# a_1359_n188# a_2703_n188# a_n2241_n100# a_2319_n188#
+ a_n849_122# a_2799_122# a_n753_n188# a_n369_n188# a_2415_122# a_n33_n100# a_735_n100#
+ a_1887_n100# a_n2193_122# a_2847_n100# a_687_122# a_n1809_122# a_303_122# a_n2673_n188#
+ a_n2289_n188# a_n1713_n188# a_n897_n100# a_n1329_n188# a_1647_122# a_831_n100# a_447_n100#
+ a_1983_n100# a_1599_n100# a_1551_n188# a_n1041_122# a_1167_n188# a_2511_n188# a_2559_n100#
+ a_2127_n188# a_n1857_n100# a_n81_122# a_15_n188# a_n2817_n100# a_n993_n100# a_2607_122#
+ a_n561_n188# a_n177_n188# a_n2385_122#
X0 a_63_n100# a_15_n188# a_n33_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n2721_n100# a_n2769_122# a_n2817_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_n2433_n100# a_n2481_n188# a_n2529_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n2241_n100# a_n2289_n188# a_n2337_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_n2145_n100# a_n2193_122# a_n2241_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_n2049_n100# a_n2097_n188# a_n2145_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n2817_n100# a_n2865_n188# a_n2909_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X7 a_n2625_n100# a_n2673_n188# a_n2721_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X8 a_n2529_n100# a_n2577_122# a_n2625_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X9 a_n2337_n100# a_n2385_122# a_n2433_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_2175_n100# a_2127_n188# a_2079_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X11 a_2271_n100# a_2223_122# a_2175_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_2463_n100# a_2415_122# a_2367_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_2751_n100# a_2703_n188# a_2655_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X14 a_2079_n100# a_2031_122# a_1983_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X15 a_2367_n100# a_2319_n188# a_2271_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X16 a_2559_n100# a_2511_n188# a_2463_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_2655_n100# a_2607_122# a_2559_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X18 a_2847_n100# a_2799_122# a_2751_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X19 a_1023_n100# a_975_n188# a_927_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X20 a_927_n100# a_879_122# a_831_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_n1761_n100# a_n1809_122# a_n1857_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X22 a_n1953_n100# a_n2001_122# a_n2049_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X23 a_n1857_n100# a_n1905_n188# a_n1953_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X24 a_n1665_n100# a_n1713_n188# a_n1761_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_n1569_n100# a_n1617_122# a_n1665_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_1215_n100# a_1167_n188# a_1119_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X27 a_1311_n100# a_1263_122# a_1215_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_1503_n100# a_1455_122# a_1407_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X29 a_1791_n100# a_1743_n188# a_1695_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X30 a_1119_n100# a_1071_122# a_1023_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_1407_n100# a_1359_n188# a_1311_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_1599_n100# a_1551_n188# a_1503_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_1695_n100# a_1647_122# a_1599_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X34 a_1887_n100# a_1839_122# a_1791_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X35 a_1983_n100# a_1935_n188# a_1887_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X36 a_n33_n100# a_n81_122# a_n129_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X37 a_351_n100# a_303_122# a_255_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X38 a_159_n100# a_111_122# a_63_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X39 a_255_n100# a_207_n188# a_159_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_447_n100# a_399_n188# a_351_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X41 a_543_n100# a_495_122# a_447_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X42 a_735_n100# a_687_122# a_639_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X43 a_831_n100# a_783_n188# a_735_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_639_n100# a_591_n188# a_543_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_n1473_n100# a_n1521_n188# a_n1569_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X46 a_n1281_n100# a_n1329_n188# a_n1377_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X47 a_n1185_n100# a_n1233_122# a_n1281_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X48 a_n993_n100# a_n1041_122# a_n1089_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X49 a_n1377_n100# a_n1425_122# a_n1473_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n1089_n100# a_n1137_n188# a_n1185_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X51 a_n321_n100# a_n369_n188# a_n417_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X52 a_n801_n100# a_n849_122# a_n897_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X53 a_n705_n100# a_n753_n188# a_n801_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X54 a_n513_n100# a_n561_n188# a_n609_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X55 a_n417_n100# a_n465_122# a_n513_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_n225_n100# a_n273_122# a_n321_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X57 a_n129_n100# a_n177_n188# a_n225_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_n897_n100# a_n945_n188# a_n993_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_n609_n100# a_n657_122# a_n705_n100# a_n3011_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_HNLS5R a_159_n100# a_n323_n274# a_n129_n100# a_n221_n100#
+ a_63_n100# a_n33_n100# a_n81_122# a_n177_n188#
X0 a_63_n100# a_n177_n188# a_n33_n100# a_n323_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_122# a_n129_n100# a_n323_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_159_n100# a_n81_122# a_63_n100# a_n323_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X3 a_n129_n100# a_n177_n188# a_n221_n100# a_n323_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
.ends

.subckt output_buffer INB INA VDD BIAS OUTB GND OUTA SUB
XXR1 VDD m1_12140_1165# SUB sky130_fd_pr__res_high_po_2p85_P79JE3
XXR2 VDD m1_12140_n1090# SUB sky130_fd_pr__res_high_po_2p85_P79JE3
XXR3 VDD OUTB SUB sky130_fd_pr__res_high_po_5p73_W59YBA
XXM1 m1_9850_15# m1_9850_15# m1_9850_15# GND GND m1_9850_15# m1_9850_15# m1_9850_15#
+ GND GND m1_9850_15# GND m1_9850_15# BIAS m1_9850_15# SUB GND GND m1_9850_15# m1_9850_15#
+ GND GND GND sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM2 m1_9850_15# m1_9850_15# m1_9850_15# GND GND m1_9850_15# m1_9850_15# m1_9850_15#
+ GND GND m1_9850_15# GND m1_9850_15# BIAS m1_9850_15# SUB GND GND m1_9850_15# m1_9850_15#
+ GND GND GND sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM3 m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15# BIAS BIAS m1_13690_15# BIAS
+ BIAS m1_13690_15# BIAS m1_13690_15# BIAS BIAS m1_13690_15# BIAS GND GND BIAS GND
+ BIAS GND GND GND BIAS GND GND BIAS m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS m1_13690_15# BIAS m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS GND BIAS GND BIAS GND BIAS GND GND GND BIAS GND GND GND BIAS m1_13690_15#
+ m1_13690_15# m1_13690_15# BIAS BIAS BIAS m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS BIAS BIAS SUB BIAS GND BIAS BIAS BIAS GND GND BIAS BIAS GND BIAS
+ BIAS GND BIAS BIAS BIAS BIAS BIAS BIAS m1_13690_15# m1_13690_15# m1_13690_15# BIAS
+ m1_13690_15# BIAS BIAS BIAS BIAS BIAS BIAS GND BIAS BIAS GND GND GND GND BIAS BIAS
+ BIAS BIAS GND BIAS GND BIAS BIAS GND m1_13690_15# BIAS BIAS BIAS BIAS sky130_fd_pr__nfet_01v8_lvt_LELFGX
XXM4 m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15# BIAS BIAS m1_13690_15# BIAS
+ BIAS m1_13690_15# BIAS m1_13690_15# BIAS BIAS m1_13690_15# BIAS GND GND BIAS GND
+ BIAS GND GND GND BIAS GND GND BIAS m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS m1_13690_15# BIAS m1_13690_15# m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS GND BIAS GND BIAS GND BIAS GND GND GND BIAS GND GND GND BIAS m1_13690_15#
+ m1_13690_15# m1_13690_15# BIAS BIAS BIAS m1_13690_15# m1_13690_15# m1_13690_15#
+ m1_13690_15# BIAS BIAS BIAS SUB BIAS GND BIAS BIAS BIAS GND GND BIAS BIAS GND BIAS
+ BIAS GND BIAS BIAS BIAS BIAS BIAS BIAS m1_13690_15# m1_13690_15# m1_13690_15# BIAS
+ m1_13690_15# BIAS BIAS BIAS BIAS BIAS BIAS GND BIAS BIAS GND GND GND GND BIAS BIAS
+ BIAS BIAS GND BIAS GND BIAS BIAS GND m1_13690_15# BIAS BIAS BIAS BIAS sky130_fd_pr__nfet_01v8_lvt_LELFGX
XXR29 VDD OUTA SUB sky130_fd_pr__res_high_po_5p73_W59YBA
XXM42 m1_9850_15# SUB m1_12140_1165# m1_9850_15# m1_12140_1165# m1_9850_15# INA INA
+ sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM43 m1_9850_15# SUB m1_12140_n1090# m1_9850_15# m1_12140_n1090# m1_9850_15# INB
+ INB sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM32 m1_13690_15# m1_13690_15# m1_13690_15# OUTA OUTA m1_13690_15# m1_13690_15# m1_13690_15#
+ OUTA OUTA m1_13690_15# OUTA m1_13690_15# m1_12140_1165# m1_13690_15# SUB OUTA OUTA
+ m1_13690_15# m1_13690_15# OUTA OUTA OUTA sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM33 m1_13690_15# m1_13690_15# m1_13690_15# OUTB OUTB m1_13690_15# m1_13690_15# m1_13690_15#
+ OUTB OUTB m1_13690_15# OUTB m1_13690_15# m1_12140_n1090# m1_13690_15# SUB OUTB OUTB
+ m1_13690_15# m1_13690_15# OUTB OUTB OUTB sky130_fd_pr__nfet_01v8_lvt_YTLFGX
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3M934 a_35_n100# a_n547_n197# a_n931_n197# a_931_n100#
+ a_547_n100# a_605_n197# a_n477_n100# a_n861_n100# a_n291_n197# a_291_n100# w_n1127_n319#
+ a_n221_n100# a_n989_n100# a_n803_n197# a_861_n197# a_n419_n197# a_477_n197# a_803_n100#
+ a_419_n100# a_n349_n100# a_n733_n100# a_n163_n197# a_163_n100# a_221_n197# a_n93_n100#
+ a_n675_n197# a_675_n100# a_733_n197# a_349_n197# a_n605_n100# a_n35_n197# a_93_n197#
X0 a_291_n100# a_221_n197# a_163_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_675_n100# a_605_n197# a_547_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X2 a_n221_n100# a_n291_n197# a_n349_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X3 a_n605_n100# a_n675_n197# a_n733_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X4 a_931_n100# a_861_n197# a_803_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_547_n100# a_477_n197# a_419_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X6 a_n93_n100# a_n163_n197# a_n221_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X7 a_163_n100# a_93_n197# a_35_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X8 a_n861_n100# a_n931_n197# a_n989_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X9 a_n477_n100# a_n547_n197# a_n605_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X10 a_419_n100# a_349_n197# a_291_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X11 a_803_n100# a_733_n197# a_675_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X12 a_35_n100# a_n35_n197# a_n93_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X13 a_n733_n100# a_n803_n197# a_n861_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X14 a_n349_n100# a_n419_n197# a_n477_n100# w_n1127_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3Z634 a_483_n100# a_1693_n197# a_541_n197# a_157_n197#
+ a_1635_n100# a_1309_n197# a_99_n100# a_n413_n100# a_n995_n197# a_n1891_n197# a_n29_n100#
+ a_n1507_n197# a_995_n100# a_1053_n197# a_669_n197# a_n925_n100# a_n1437_n100# a_n1821_n100#
+ w_n2087_n319# a_n355_n197# a_n1251_n197# a_413_n197# a_1891_n100# a_355_n100# a_n1181_n100#
+ a_1565_n197# a_1507_n100# a_n285_n100# a_29_n197# a_n1949_n100# a_n1763_n197# a_n867_n197#
+ a_n1379_n197# a_1251_n100# a_867_n100# a_925_n197# a_n797_n100# a_n1693_n100# a_n1309_n100#
+ a_n227_n197# a_n611_n197# a_n1123_n197# a_285_n197# a_1763_n100# a_1379_n100# a_611_n100#
+ a_227_n100# a_1821_n197# a_1437_n197# a_n157_n100# a_n541_n100# a_n1053_n100# a_n1635_n197#
+ a_n739_n197# a_1181_n197# a_797_n197# a_739_n100# a_1123_n100# a_n1565_n100# a_n669_n100#
+ a_n483_n197# a_n99_n197#
X0 a_483_n100# a_413_n197# a_355_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n1181_n100# a_n1251_n197# a_n1309_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X2 a_n1565_n100# a_n1635_n197# a_n1693_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X3 a_n413_n100# a_n483_n197# a_n541_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X4 a_n797_n100# a_n867_n197# a_n925_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X5 a_355_n100# a_285_n197# a_227_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X6 a_739_n100# a_669_n197# a_611_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X7 a_n1821_n100# a_n1891_n197# a_n1949_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X8 a_1123_n100# a_1053_n197# a_995_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X9 a_1507_n100# a_1437_n197# a_1379_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X10 a_1891_n100# a_1821_n197# a_1763_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X11 a_99_n100# a_29_n197# a_n29_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X12 a_1763_n100# a_1693_n197# a_1635_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X13 a_n1053_n100# a_n1123_n197# a_n1181_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X14 a_n1437_n100# a_n1507_n197# a_n1565_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X15 a_n285_n100# a_n355_n197# a_n413_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X16 a_n669_n100# a_n739_n197# a_n797_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X17 a_611_n100# a_541_n197# a_483_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X18 a_227_n100# a_157_n197# a_99_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X19 a_995_n100# a_925_n197# a_867_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X20 a_n1693_n100# a_n1763_n197# a_n1821_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X21 a_n1309_n100# a_n1379_n197# a_n1437_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X22 a_n925_n100# a_n995_n197# a_n1053_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X23 a_1379_n100# a_1309_n197# a_1251_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X24 a_867_n100# a_797_n197# a_739_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X25 a_1251_n100# a_1181_n197# a_1123_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X26 a_1635_n100# a_1565_n197# a_1507_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X27 a_n541_n100# a_n611_n197# a_n669_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X28 a_n157_n100# a_n227_n197# a_n285_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X29 a_n29_n100# a_n99_n197# a_n157_n100# w_n2087_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_9DHFGX a_159_n100# a_111_n188# a_15_122# a_n273_n188#
+ a_255_n100# a_n611_n274# a_351_n100# a_n417_n100# a_207_122# a_n129_n100# a_n81_n188#
+ a_63_n100# a_n177_122# a_n225_n100# a_n321_n100# a_n369_122# a_n33_n100# a_n509_n100#
+ a_303_n188# a_n465_n188# a_447_n100# a_399_122#
X0 a_63_n100# a_15_122# a_n33_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_n188# a_n129_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_351_n100# a_303_n188# a_255_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_159_n100# a_111_n188# a_63_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_255_n100# a_207_122# a_159_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_447_n100# a_399_122# a_351_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_n321_n100# a_n369_122# a_n417_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X7 a_n417_n100# a_n465_n188# a_n509_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X8 a_n225_n100# a_n273_n188# a_n321_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X9 a_n129_n100# a_n177_122# a_n225_n100# a_n611_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_MM89SS a_n285_n1572# a_n415_n1702# a_n285_1140#
X0 a_n285_n1572# a_n285_1140# a_n415_n1702# sky130_fd_pr__res_high_po_2p85 l=1.14e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4 a_483_n100# a_541_n197# a_157_n197# a_99_n100#
+ a_n413_n100# a_n29_n100# a_n355_n197# a_413_n197# a_355_n100# a_n285_n100# a_29_n197#
+ w_n807_n319# a_n227_n197# a_n611_n197# a_285_n197# a_611_n100# a_227_n100# a_n157_n100#
+ a_n541_n100# a_n669_n100# a_n483_n197# a_n99_n197#
X0 a_483_n100# a_413_n197# a_355_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_n413_n100# a_n483_n197# a_n541_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X2 a_355_n100# a_285_n197# a_227_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X3 a_99_n100# a_29_n197# a_n29_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X4 a_n285_n100# a_n355_n197# a_n413_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X5 a_611_n100# a_541_n197# a_483_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X6 a_227_n100# a_157_n197# a_99_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
X7 a_n541_n100# a_n611_n197# a_n669_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X8 a_n157_n100# a_n227_n197# a_n285_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=350000u
X9 a_n29_n100# a_n99_n197# a_n157_n100# w_n807_n319# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt bias_calc AMP VCTRL PSUB BIASOUT VOP VDD BIAS2V GND SUB
XXM36 m1_17310_5240# BIAS2V BIAS2V VDD m1_17310_5240# BIAS2V m1_17310_5240# VDD BIAS2V
+ m1_17310_5240# PSUB m1_17310_5240# m1_17310_5240# BIAS2V BIAS2V BIAS2V BIAS2V m1_17310_5240#
+ VDD VDD m1_17310_5240# BIAS2V VDD BIAS2V VDD BIAS2V VDD BIAS2V BIAS2V VDD BIAS2V
+ BIAS2V sky130_fd_pr__pfet_01v8_lvt_D3M934
XXM37 m1_17310_5240# VCTRL VCTRL VCTRL m1_17860_4190# VCTRL m1_17860_4190# m1_17860_4190#
+ VCTRL VCTRL m1_17310_5240# VCTRL m1_17310_5240# VCTRL VCTRL m1_17860_4190# m1_17860_4190#
+ m1_17310_5240# PSUB VCTRL VCTRL VCTRL m1_17860_4190# m1_17860_4190# m1_17860_4190#
+ VCTRL m1_17310_5240# m1_17310_5240# VCTRL m1_17860_4190# VCTRL VCTRL VCTRL m1_17310_5240#
+ m1_17860_4190# VCTRL m1_17310_5240# m1_17860_4190# m1_17310_5240# VCTRL VCTRL VCTRL
+ VCTRL m1_17310_5240# m1_17860_4190# m1_17860_4190# m1_17310_5240# VCTRL VCTRL m1_17860_4190#
+ m1_17310_5240# m1_17310_5240# VCTRL VCTRL VCTRL VCTRL m1_17310_5240# m1_17860_4190#
+ m1_17310_5240# m1_17860_4190# VCTRL VCTRL sky130_fd_pr__pfet_01v8_lvt_D3Z634
XXM38 m1_17310_5240# m1_18270_400# m1_18270_400# m1_18270_400# BIASOUT m1_18270_400#
+ BIASOUT BIASOUT m1_18270_400# m1_18270_400# m1_17310_5240# m1_18270_400# m1_17310_5240#
+ m1_18270_400# m1_18270_400# BIASOUT BIASOUT m1_17310_5240# PSUB m1_18270_400# m1_18270_400#
+ m1_18270_400# BIASOUT BIASOUT BIASOUT m1_18270_400# m1_17310_5240# m1_17310_5240#
+ m1_18270_400# BIASOUT m1_18270_400# m1_18270_400# m1_18270_400# m1_17310_5240# BIASOUT
+ m1_18270_400# m1_17310_5240# BIASOUT m1_17310_5240# m1_18270_400# m1_18270_400#
+ m1_18270_400# m1_18270_400# m1_17310_5240# BIASOUT BIASOUT m1_17310_5240# m1_18270_400#
+ m1_18270_400# BIASOUT m1_17310_5240# m1_17310_5240# m1_18270_400# m1_18270_400#
+ m1_18270_400# m1_18270_400# m1_17310_5240# BIASOUT m1_17310_5240# BIASOUT m1_18270_400#
+ m1_18270_400# sky130_fd_pr__pfet_01v8_lvt_D3Z634
XXM39 m1_17860_4190# m1_17860_4190# m1_17860_4190# m1_17860_4190# GND SUB m1_17860_4190#
+ m1_17860_4190# m1_17860_4190# GND m1_17860_4190# GND m1_17860_4190# m1_17860_4190#
+ GND m1_17860_4190# m1_17860_4190# GND m1_17860_4190# m1_17860_4190# GND m1_17860_4190#
+ sky130_fd_pr__nfet_01v8_lvt_9DHFGX
XXM29 VDD BIAS2V BIAS2V m1_20160_2025# VDD BIAS2V VDD m1_20160_2025# BIAS2V VDD PSUB
+ VDD VDD BIAS2V BIAS2V BIAS2V BIAS2V VDD m1_20160_2025# m1_20160_2025# VDD BIAS2V
+ m1_20160_2025# BIAS2V m1_20160_2025# BIAS2V m1_20160_2025# BIAS2V BIAS2V m1_20160_2025#
+ BIAS2V BIAS2V sky130_fd_pr__pfet_01v8_lvt_D3M934
XXR20 m1_18270_400# SUB GND sky130_fd_pr__res_high_po_2p85_MM89SS
XXM1 m1_20160_2025# BIAS2V BIAS2V VDD m1_20160_2025# BIAS2V m1_20160_2025# VDD BIAS2V
+ m1_20160_2025# PSUB m1_20160_2025# m1_20160_2025# BIAS2V BIAS2V BIAS2V BIAS2V m1_20160_2025#
+ VDD VDD m1_20160_2025# BIAS2V VDD BIAS2V VDD BIAS2V VDD BIAS2V BIAS2V VDD BIAS2V
+ BIAS2V sky130_fd_pr__pfet_01v8_lvt_D3M934
XXM2 m1_17310_5240# BIAS2V BIAS2V VDD m1_17310_5240# BIAS2V m1_17310_5240# VDD BIAS2V
+ m1_17310_5240# PSUB m1_17310_5240# m1_17310_5240# BIAS2V BIAS2V BIAS2V BIAS2V m1_17310_5240#
+ VDD VDD m1_17310_5240# BIAS2V VDD BIAS2V VDD BIAS2V VDD BIAS2V BIAS2V VDD BIAS2V
+ BIAS2V sky130_fd_pr__pfet_01v8_lvt_D3M934
XXM3 m1_17310_5240# BIAS2V BIAS2V VDD m1_17310_5240# BIAS2V m1_17310_5240# VDD BIAS2V
+ m1_17310_5240# PSUB m1_17310_5240# m1_17310_5240# BIAS2V BIAS2V BIAS2V BIAS2V m1_17310_5240#
+ VDD VDD m1_17310_5240# BIAS2V VDD BIAS2V VDD BIAS2V VDD BIAS2V BIAS2V VDD BIAS2V
+ BIAS2V sky130_fd_pr__pfet_01v8_lvt_D3M934
XXR19 GND m1_19235_6325# SUB sky130_fd_pr__res_high_po_2p85_P79JE3
XXM40 BIASOUT m1_17860_4190# m1_17860_4190# m1_17860_4190# GND SUB BIASOUT BIASOUT
+ m1_17860_4190# GND m1_17860_4190# GND m1_17860_4190# BIASOUT GND m1_17860_4190#
+ BIASOUT GND m1_17860_4190# m1_17860_4190# GND m1_17860_4190# sky130_fd_pr__nfet_01v8_lvt_9DHFGX
XXM30 m1_18270_400# VOP VOP m1_20160_2025# m1_20160_2025# m1_18270_400# VOP VOP m1_20160_2025#
+ m1_18270_400# VOP PSUB VOP VOP VOP m1_20160_2025# m1_18270_400# m1_20160_2025# m1_18270_400#
+ m1_20160_2025# VOP VOP sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4
XXM31 m1_19235_6325# AMP AMP m1_20160_2025# m1_20160_2025# m1_19235_6325# AMP AMP
+ m1_20160_2025# m1_19235_6325# AMP PSUB AMP AMP AMP m1_20160_2025# m1_19235_6325#
+ m1_20160_2025# m1_19235_6325# m1_20160_2025# AMP AMP sky130_fd_pr__pfet_01v8_lvt_D3ZSZ4
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_75KH85 a_n93_n64# a_n35_n161# a_93_n161# w_n359_n284#
+ a_35_n64# a_n163_n161# a_n221_n64# a_163_n64#
X0 a_n93_n64# a_n163_n161# a_n221_n64# w_n359_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X1 a_163_n64# a_93_n161# a_35_n64# w_n359_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=350000u
X2 a_35_n64# a_n35_n161# a_n93_n64# w_n359_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=350000u
.ends

.subckt core_osc_amp INB INA VDD BIAS GND OUTB OUTA SUB
XXM1 m1_3550_1144# m1_3550_1144# m1_3550_1144# GND GND m1_3550_1144# m1_3550_1144#
+ m1_3550_1144# GND GND m1_3550_1144# GND m1_3550_1144# BIAS m1_3550_1144# SUB GND
+ GND m1_3550_1144# m1_3550_1144# GND GND GND sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXM2 OUTA SUB m1_3550_1144# OUTA m1_3550_1144# OUTA INA INA sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM3 OUTB SUB m1_3550_1144# OUTB m1_3550_1144# OUTB INB INB sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXR16 VDD OUTA SUB sky130_fd_pr__res_high_po_2p85_P79JE3
XXM4 m1_3550_1144# m1_3550_1144# m1_3550_1144# GND GND m1_3550_1144# m1_3550_1144#
+ m1_3550_1144# GND GND m1_3550_1144# GND m1_3550_1144# BIAS m1_3550_1144# SUB GND
+ GND m1_3550_1144# m1_3550_1144# GND GND GND sky130_fd_pr__nfet_01v8_lvt_YTLFGX
XXR17 VDD OUTB SUB sky130_fd_pr__res_high_po_2p85_P79JE3
.ends

.subckt core_osc VDD GND S1B S1A S3A S3B S4B S4A BIAS S2B S2A SUB
XX4 S3B S3A VDD BIAS GND S4B S4A SUB core_osc_amp
XX1 S4A S4B VDD BIAS GND S1B S1A SUB core_osc_amp
XX2 S1B S1A VDD BIAS GND S2B S2A SUB core_osc_amp
XX3 S2B S2A VDD BIAS GND S3B S3A SUB core_osc_amp
.ends

.subckt sky130_fd_pr__res_high_po_5p73_YZEQ6M a_n573_n3472# a_n703_n3602# a_n573_3040#
X0 a_n573_n3472# a_n573_3040# a_n703_n3602# sky130_fd_pr__res_high_po_5p73 l=3.04e+07u
.ends

.subckt buffer_amp INB INA VDD BIAS OUTB GND OUTA SUB
XXR1 OUTB SUB VDD sky130_fd_pr__res_high_po_5p73_YZEQ6M
XXR2 OUTA SUB VDD sky130_fd_pr__res_high_po_5p73_YZEQ6M
XXM1 m1_6810_1630# BIAS BIAS BIAS GND SUB m1_6810_1630# m1_6810_1630# BIAS GND BIAS
+ GND BIAS m1_6810_1630# GND BIAS m1_6810_1630# GND BIAS BIAS GND BIAS sky130_fd_pr__nfet_01v8_lvt_9DHFGX
XXM2 m1_6810_1630# INB OUTB SUB sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM3 m1_6810_1630# INA OUTA SUB sky130_fd_pr__nfet_01v8_lvt_648S5X
XXM4 m1_6810_1630# BIAS BIAS BIAS GND SUB m1_6810_1630# m1_6810_1630# BIAS GND BIAS
+ GND BIAS m1_6810_1630# GND BIAS m1_6810_1630# GND BIAS BIAS GND BIAS sky130_fd_pr__nfet_01v8_lvt_9DHFGX
.ends

.subckt sky130_fd_pr__res_high_po_2p85_MXEQGY a_n285_4200# a_n285_n4632# a_n415_n4762#
X0 a_n285_n4632# a_n285_4200# a_n415_n4762# sky130_fd_pr__res_high_po_2p85 l=4.2e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_4RCNTW c1_n2050_n3000# m3_n2150_n3100#
X0 c1_n2050_n3000# m3_n2150_n3100# sky130_fd_pr__cap_mim_m3_1 l=3e+07u w=2e+07u
.ends

.subckt amp_dec AMP IN4 IN3 IN2 IN1 VDD GND SUB
XXM25 AMP SUB VDD AMP VDD AMP IN3 IN3 sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM26 AMP SUB VDD AMP VDD AMP IN4 IN4 sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM27 AMP SUB VDD AMP VDD AMP IN2 IN2 sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXM28 AMP SUB VDD AMP VDD AMP IN1 IN1 sky130_fd_pr__nfet_01v8_lvt_HNLS5R
XXR18 AMP GND SUB sky130_fd_pr__res_high_po_2p85_MXEQGY
XXC1 AMP GND sky130_fd_pr__cap_mim_m3_1_4RCNTW
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_6BNFGK a_543_n100# a_159_n100# a_n273_122# a_255_n100#
+ a_351_n100# a_n417_n100# a_n465_122# a_n129_n100# a_n513_n100# a_399_n188# a_63_n100#
+ a_n225_n100# a_495_122# a_111_122# a_n321_n100# a_207_n188# a_n369_n188# a_n33_n100#
+ a_n707_n274# a_303_122# a_n605_n100# a_447_n100# a_15_n188# a_n81_122# a_n177_n188#
+ a_n561_n188#
X0 a_63_n100# a_15_n188# a_n33_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n33_n100# a_n81_122# a_n129_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_351_n100# a_303_122# a_255_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_159_n100# a_111_122# a_63_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_255_n100# a_207_n188# a_159_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X5 a_447_n100# a_399_n188# a_351_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X6 a_543_n100# a_495_122# a_447_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_n321_n100# a_n369_n188# a_n417_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X8 a_n513_n100# a_n561_n188# a_n605_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X9 a_n417_n100# a_n465_122# a_n513_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n225_n100# a_n273_122# a_n321_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_n129_n100# a_n177_n188# a_n225_n100# a_n707_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt vop_dec VOP VDD IN GND SUB
XXR21 VOP GND SUB sky130_fd_pr__res_high_po_2p85_MXEQGY
XXC2 IN GND sky130_fd_pr__cap_mim_m3_1_4RCNTW
XXM41 VDD VDD IN VOP VDD VDD IN VOP VOP IN VOP VDD IN IN VOP IN IN VDD SUB IN VDD
+ VOP IN IN IN IN sky130_fd_pr__nfet_01v8_lvt_6BNFGK
.ends

.subckt buffer_amp_vop I1A I1B AMP I3B I3A I4B I4A OUT0 I2B I2A VOP OUT180 BIAS GND
+ VDD SUB
XX4 I4B I4A VDD BIAS X6/IN GND X6/IN SUB buffer_amp
XX5 AMP OUT270 OUT90 OUT0 OUT180 VDD GND SUB amp_dec
XX6 VOP VDD X6/IN GND SUB vop_dec
XX1 I1B I1A VDD BIAS OUT180 GND OUT0 SUB buffer_amp
XX2 I2B I2A VDD BIAS X6/IN GND X6/IN SUB buffer_amp
XX3 I3B I3A VDD BIAS OUT270 GND OUT90 SUB buffer_amp
.ends

.subckt VCO bias_calc_0/BIAS2V CTRL5 CTRL4 bias_calc_0/VCTRL CTRL3 VDD output_buffer_0/OUTB
+ CTRL2 output_buffer_0/OUTA CTRL1 GND
XX4 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X4/IN GND cap_bank
XX5 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X5/IN GND cap_bank
XX6 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X6/IN GND cap_bank
Xoutput_buffer_0 X3/OUT180 X3/OUT0 VDD X3/BIAS output_buffer_0/OUTB GND output_buffer_0/OUTA
+ GND output_buffer
XX10 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X3/I4B GND cap_bank
XX7 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X7/IN GND cap_bank
XX8 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X8/IN GND cap_bank
XX11 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X3/I4A GND cap_bank
XX9 CTRL5 CTRL4 CTRL2 CTRL3 CTRL1 X9/IN GND cap_bank
Xbias_calc_0 X3/AMP bias_calc_0/VCTRL VDD X3/BIAS X3/VOP VDD bias_calc_0/BIAS2V GND
+ GND bias_calc
Xsky130_fd_pr__pfet_01v8_lvt_75KH85_0 VDD bias_calc_0/BIAS2V bias_calc_0/BIAS2V VDD
+ bias_calc_0/BIAS2V bias_calc_0/BIAS2V bias_calc_0/BIAS2V VDD sky130_fd_pr__pfet_01v8_lvt_75KH85
XX1 VDD GND X4/IN X5/IN X9/IN X8/IN X3/I4B X3/I4A X3/BIAS X6/IN X7/IN GND core_osc
XX3 X5/IN X4/IN X3/AMP X8/IN X9/IN X3/I4B X3/I4A X3/OUT0 X6/IN X7/IN X3/VOP X3/OUT180
+ X3/BIAS GND VDD GND buffer_amp_vop
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_M9466H a_100_n200# a_n158_n200# a_n100_n288# a_n260_n374#
X0 a_100_n200# a_n100_n288# a_n158_n200# a_n260_n374# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
.ends

.subckt TX_line INB OUTA VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_M9466H_0 VSUBS VSUBS VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt_M9466H
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_UZMRKM a_669_10600# a_n3057_n11032# a_n1815_n11032#
+ a_n3057_10600# a_n1815_10600# a_n3187_n11162# a_669_n11032# a_n573_10600# a_n573_n11032#
+ a_1911_n11032# a_1911_10600#
X0 a_n3057_n11032# a_n3057_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X1 a_n573_n11032# a_n573_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X2 a_n1815_n11032# a_n1815_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X3 a_669_n11032# a_669_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
X4 a_1911_n11032# a_1911_10600# a_n3187_n11162# sky130_fd_pr__res_xhigh_po_5p73 l=1.06e+08u
.ends

.subckt XM_Rref sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_1911_n11032# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_n3057_10600#
+ VSUBS
Xsky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0 m1_3616_20636# m1_n110_n995# m1_n110_n995#
+ sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_n3057_10600# m1_1132_20636# VSUBS m1_2374_n995#
+ m1_1132_20636# m1_2374_n995# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM_0/a_1911_n11032#
+ m1_3616_20636# sky130_fd_pr__res_xhigh_po_5p73_UZMRKM
.ends

.subckt sky130_fd_pr__res_high_po_1p41_S8KB58 a_n141_n4671# a_n141_4239# a_n271_n4801#
X0 a_n141_n4671# a_n141_4239# a_n271_n4801# sky130_fd_pr__res_high_po_1p41 l=4.239e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_TSNZVH a_50_n364# w_n246_n584# a_n108_n364# a_n50_n461#
X0 a_50_n364# a_n50_n461# a_n108_n364# w_n246_n584# sky130_fd_pr__pfet_01v8 ad=1.16e+12p pd=8.58e+06u as=1.16e+12p ps=8.58e+06u w=4e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_Y5UG24 a_n108_n181# a_n50_n207# a_n210_n293# a_50_n181#
X0 a_50_n181# a_n50_n207# a_n108_n181# a_n210_n293# sky130_fd_pr__nfet_01v8 ad=4.35e+11p pd=3.58e+06u as=4.35e+11p ps=3.58e+06u w=1.5e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_high_po_1p41_2TBR6S a_n141_n2032# a_n141_1600# a_n271_n2162#
X0 a_n141_n2032# a_n141_1600# a_n271_n2162# sky130_fd_pr__res_high_po_1p41 l=1.6e+07u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_Y9W37A m3_n2450_n680# c1_n2350_n580#
X0 c1_n2350_n580# m3_n2450_n680# sky130_fd_pr__cap_mim_m3_1 l=5.8e+06u w=2.3e+07u
.ends

.subckt XM_pdn sky130_fd_pr__cap_mim_m3_1_Y9W37A_0/c1_n2350_n580# sky130_fd_pr__nfet_01v8_Y5UG24_2/a_n108_n181#
+ m1_160_n220# li_97_967# sky130_fd_pr__nfet_01v8_Y5UG24_2/a_50_n181# VSUBS
Xsky130_fd_pr__pfet_01v8_TSNZVH_0 m1_280_n320# li_97_967# li_97_967# m1_160_n220#
+ sky130_fd_pr__pfet_01v8_TSNZVH
Xsky130_fd_pr__pfet_01v8_TSNZVH_1 m1_660_n320# li_97_967# li_97_967# m1_280_n320#
+ sky130_fd_pr__pfet_01v8_TSNZVH
Xsky130_fd_pr__nfet_01v8_Y5UG24_0 VSUBS m1_160_n220# VSUBS m1_280_n320# sky130_fd_pr__nfet_01v8_Y5UG24
Xsky130_fd_pr__nfet_01v8_Y5UG24_1 VSUBS m1_280_n320# VSUBS m1_660_n320# sky130_fd_pr__nfet_01v8_Y5UG24
Xsky130_fd_pr__nfet_01v8_Y5UG24_2 sky130_fd_pr__nfet_01v8_Y5UG24_2/a_n108_n181# m1_910_n240#
+ VSUBS sky130_fd_pr__nfet_01v8_Y5UG24_2/a_50_n181# sky130_fd_pr__nfet_01v8_Y5UG24
Xsky130_fd_pr__res_high_po_1p41_2TBR6S_0 m1_660_n320# m1_910_n240# VSUBS sky130_fd_pr__res_high_po_1p41_2TBR6S
Xsky130_fd_pr__cap_mim_m3_1_Y9W37A_0 m1_910_n240# sky130_fd_pr__cap_mim_m3_1_Y9W37A_0/c1_n2350_n580#
+ sky130_fd_pr__cap_mim_m3_1_Y9W37A
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_Q24T46 a_n416_n136# a_n616_n162# w_n812_n284#
+ a_358_n136# a_158_n162# a_100_n136# a_n674_n136# a_n158_n136# a_n358_n162# a_616_n136#
+ a_416_n162# a_n100_n162#
X0 a_358_n136# a_158_n162# a_100_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_616_n136# a_416_n162# a_358_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X2 a_100_n136# a_n100_n162# a_n158_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_n416_n136# a_n616_n162# a_n674_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_n158_n136# a_n358_n162# a_n416_n136# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MUVY4U a_n616_n161# a_358_n64# a_n674_n64# a_n158_n64#
+ w_n812_n284# a_158_n161# a_n358_n161# a_416_n161# a_n100_n161# a_616_n64# a_100_n64#
+ a_n416_n64#
X0 a_100_n64# a_n100_n161# a_n158_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_616_n64# a_416_n161# a_358_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_358_n64# a_158_n161# a_100_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X3 a_n416_n64# a_n616_n161# a_n674_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_n158_n64# a_n358_n161# a_n416_n64# w_n812_n284# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt XM_current_gate m1_30_n420# m1_94_n180# li_818_316# m1_30_260#
Xsky130_fd_pr__pfet_01v8_lvt_Q24T46_0 li_818_316# m1_94_n180# li_818_316# m1_30_n420#
+ m1_94_n180# li_818_316# m1_30_n420# m1_30_260# m1_94_n180# li_818_316# m1_94_n180#
+ m1_94_n180# sky130_fd_pr__pfet_01v8_lvt_Q24T46
Xsky130_fd_pr__pfet_01v8_lvt_MUVY4U_0 m1_94_n180# m1_30_260# m1_30_260# m1_30_n420#
+ li_818_316# m1_94_n180# m1_94_n180# m1_94_n180# m1_94_n180# li_818_316# li_818_316#
+ li_818_316# sky130_fd_pr__pfet_01v8_lvt_MUVY4U
.ends

.subckt XM_current_gate_with_dummy XM_current_gate_6/m1_30_n420# XM_current_gate_2/m1_94_n180#
+ XM_current_gate_8/m1_30_260# XM_current_gate_5/m1_94_n180# XM_current_gate_1/m1_94_n180#
+ XM_current_gate_8/m1_94_n180# XM_current_gate_3/m1_94_n180# XM_current_gate_1/m1_30_260#
+ XM_current_gate_6/m1_94_n180# XM_current_gate_7/m1_30_n420# XM_current_gate_5/m1_30_n420#
+ XM_current_gate_0/m1_30_n420# XM_current_gate_2/m1_30_260# XM_current_gate_8/m1_30_n420#
+ XM_current_gate_2/m1_30_n420# XM_current_gate_4/m1_94_n180# XM_current_gate_5/m1_30_260#
+ XM_current_gate_0/m1_94_n180# XM_current_gate_4/m1_30_260# XM_current_gate_7/m1_30_260#
+ XM_current_gate_3/m1_30_n420# XM_current_gate_8/li_818_316# XM_current_gate_4/m1_30_n420#
+ XM_current_gate_1/m1_30_n420# XM_current_gate_0/m1_30_260# XM_current_gate_3/m1_30_260#
+ XM_current_gate_6/m1_30_260# XM_current_gate_7/m1_94_n180#
XXM_current_gate_0 XM_current_gate_0/m1_30_n420# XM_current_gate_0/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_0/m1_30_260# XM_current_gate
XXM_current_gate_1 XM_current_gate_1/m1_30_n420# XM_current_gate_1/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_1/m1_30_260# XM_current_gate
XXM_current_gate_2 XM_current_gate_2/m1_30_n420# XM_current_gate_2/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_2/m1_30_260# XM_current_gate
XXM_current_gate_3 XM_current_gate_3/m1_30_n420# XM_current_gate_3/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_3/m1_30_260# XM_current_gate
XXM_current_gate_4 XM_current_gate_4/m1_30_n420# XM_current_gate_4/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_4/m1_30_260# XM_current_gate
XXM_current_gate_5 XM_current_gate_5/m1_30_n420# XM_current_gate_5/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_5/m1_30_260# XM_current_gate
XXM_current_gate_6 XM_current_gate_6/m1_30_n420# XM_current_gate_6/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_6/m1_30_260# XM_current_gate
XXM_current_gate_7 XM_current_gate_7/m1_30_n420# XM_current_gate_7/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_7/m1_30_260# XM_current_gate
XXM_current_gate_8 XM_current_gate_8/m1_30_n420# XM_current_gate_8/m1_94_n180# XM_current_gate_8/li_818_316#
+ XM_current_gate_8/m1_30_260# XM_current_gate
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_8URDWJ a_1003_n795# a_745_300# a_803_n892# a_229_1030#
+ a_545_933# w_n1097_n1260# w_n1097_n165# a_229_300# a_1003_n65# a_n287_n430# a_287_203#
+ a_1003_665# a_n1061_n430# a_n1061_300# a_n29_n795# a_n545_1030# a_287_n1257# a_487_n795#
+ a_545_568# a_n545_300# a_745_n430# a_n229_n892# a_n1061_n1160# a_n1003_n892# a_29_933#
+ a_n1003_933# a_287_n892# a_n745_203# a_1003_1030# a_29_n527# a_n803_n65# a_n803_665#
+ a_n803_n795# a_n487_n162# a_n229_203# a_487_300# a_n745_n527# w_n1097_n895# a_29_568#
+ a_n1003_568# a_287_933# a_n29_300# a_545_n1257# a_545_n162# a_n487_n1257# a_29_n1257#
+ a_745_n65# a_803_n527# a_n29_1030# a_745_665# a_229_n430# a_487_1030# a_487_n1160#
+ w_n1097_200# a_229_n65# a_229_665# a_n287_n795# a_n287_n1160# a_n287_300# a_287_568#
+ a_n1061_n795# a_n545_n430# a_803_203# a_n1061_n65# a_n745_933# a_n1061_665# a_n229_n527#
+ a_n487_203# a_n803_1030# a_n545_n65# a_n1003_n527# a_n487_n892# a_n229_933# a_n545_665#
+ a_287_n527# a_745_n795# a_1003_n430# a_n1003_n1257# a_803_n1257# a_n745_n1257# a_545_n892#
+ a_n745_568# a_29_n162# a_745_n1160# a_487_n65# w_n1097_930# a_n229_568# a_487_665#
+ a_n545_n1160# a_1003_300# a_n745_n162# a_1003_n1160# a_n287_1030# a_n29_n65# a_n1061_1030#
+ a_n29_665# a_n29_n430# a_803_933# a_487_n430# a_803_n162# a_229_n795# a_545_203#
+ a_n487_933# w_n1097_565# a_745_1030# a_n287_n65# a_n287_665# a_n545_n795# a_803_568#
+ a_n803_300# a_n229_n1257# a_n29_n1160# a_n803_n430# a_29_n892# a_n487_n527# a_n487_568#
+ a_n229_n162# a_n803_n1160# w_n1097_n530# a_229_n1160# a_n1003_n162# a_n1003_203#
+ a_29_203# a_287_n162# a_n745_n892# a_545_n527#
X0 a_n545_n795# a_n745_n892# a_n803_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_n803_n795# a_n1003_n892# a_n1061_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_n287_n795# a_n487_n892# a_n545_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X3 a_n287_n65# a_n487_n162# a_n545_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_1003_n430# a_803_n527# a_745_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X5 a_n803_665# a_n1003_568# a_n1061_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X6 a_745_665# a_545_568# a_487_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X7 a_745_n430# a_545_n527# a_487_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X8 a_n29_665# a_n229_568# a_n287_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X9 a_487_n430# a_287_n527# a_229_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X10 a_n803_300# a_n1003_203# a_n1061_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X11 a_745_300# a_545_203# a_487_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X12 a_229_665# a_29_568# a_n29_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X13 a_n29_300# a_n229_203# a_n287_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X14 a_229_300# a_29_203# a_n29_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X15 a_487_n1160# a_287_n1257# a_229_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X16 a_n29_1030# a_n229_933# a_n287_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X17 a_229_1030# a_29_933# a_n29_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X18 a_1003_n65# a_803_n162# a_745_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X19 a_745_n795# a_545_n892# a_487_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X20 a_1003_n795# a_803_n892# a_745_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X21 a_487_665# a_287_568# a_229_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X22 a_487_n795# a_287_n892# a_229_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X23 a_n287_n1160# a_n487_n1257# a_n545_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X24 a_n545_665# a_n745_568# a_n803_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X25 a_487_300# a_287_203# a_229_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X26 a_n29_n1160# a_n229_n1257# a_n287_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X27 a_n545_300# a_n745_203# a_n803_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X28 a_n545_1030# a_n745_933# a_n803_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X29 a_n803_1030# a_n1003_933# a_n1061_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X30 a_n287_1030# a_n487_933# a_n545_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X31 a_n803_n65# a_n1003_n162# a_n1061_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X32 a_745_n65# a_545_n162# a_487_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X33 a_229_n430# a_29_n527# a_n29_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X34 a_n29_n65# a_n229_n162# a_n287_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X35 a_n29_n430# a_n229_n527# a_n287_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X36 a_745_n1160# a_545_n1257# a_487_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X37 a_n287_665# a_n487_568# a_n545_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X38 a_229_n65# a_29_n162# a_n29_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X39 a_n545_n1160# a_n745_n1257# a_n803_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X40 a_229_n1160# a_29_n1257# a_n29_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X41 a_n287_300# a_n487_203# a_n545_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X42 a_487_n65# a_287_n162# a_229_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X43 a_n545_n430# a_n745_n527# a_n803_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X44 a_n287_n430# a_n487_n527# a_n545_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X45 a_n29_n795# a_n229_n892# a_n287_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X46 a_229_n795# a_29_n892# a_n29_n795# w_n1097_n895# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X47 a_745_1030# a_545_933# a_487_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X48 a_1003_1030# a_803_933# a_745_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X49 a_n803_n430# a_n1003_n527# a_n1061_n430# w_n1097_n530# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X50 a_487_1030# a_287_933# a_229_1030# w_n1097_930# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X51 a_n545_n65# a_n745_n162# a_n803_n65# w_n1097_n165# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X52 a_1003_n1160# a_803_n1257# a_745_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X53 a_1003_665# a_803_568# a_745_665# w_n1097_565# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X54 a_1003_300# a_803_203# a_745_300# w_n1097_200# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X55 a_n803_n1160# a_n1003_n1257# a_n1061_n1160# w_n1097_n1260# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
.ends

.subckt XM_feedbackmir m1_30_180# B m1_290_100# m1_290_460# m1_98_12#
Xsky130_fd_pr__pfet_01v8_lvt_8URDWJ_0 m1_30_180# m1_290_460# m1_98_12# m1_290_100#
+ m1_98_12# B B m1_290_100# m1_30_180# m1_290_460# m1_98_12# m1_30_180# m1_30_180#
+ m1_30_180# m1_30_180# m1_30_180# m1_98_12# m1_30_180# m1_98_12# m1_30_180# m1_290_460#
+ m1_98_12# m1_30_180# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_30_180#
+ m1_98_12# m1_290_460# m1_290_460# m1_290_460# m1_98_12# m1_98_12# m1_30_180# m1_98_12#
+ B m1_98_12# m1_98_12# m1_98_12# m1_30_180# m1_98_12# m1_98_12# m1_98_12# m1_98_12#
+ m1_290_100# m1_98_12# m1_30_180# m1_290_100# m1_290_100# m1_30_180# m1_30_180# B
+ m1_290_460# m1_290_460# m1_290_100# m1_290_460# m1_290_460# m1_98_12# m1_30_180#
+ m1_30_180# m1_98_12# m1_30_180# m1_98_12# m1_30_180# m1_98_12# m1_98_12# m1_290_100#
+ m1_30_180# m1_98_12# m1_98_12# m1_98_12# m1_30_180# m1_98_12# m1_290_100# m1_30_180#
+ m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_290_460# m1_30_180#
+ B m1_98_12# m1_30_180# m1_30_180# m1_30_180# m1_98_12# m1_30_180# m1_290_460# m1_30_180#
+ m1_30_180# m1_30_180# m1_30_180# m1_98_12# m1_30_180# m1_98_12# m1_290_460# m1_98_12#
+ m1_98_12# B m1_290_460# m1_290_100# m1_290_100# m1_30_180# m1_98_12# m1_290_100#
+ m1_98_12# m1_30_180# m1_290_100# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_290_100#
+ B m1_290_100# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_98_12# m1_98_12# sky130_fd_pr__pfet_01v8_lvt_8URDWJ
.ends

.subckt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 Emitter Collector Base m=1
X0 Collector Base Emitter sky130_fd_pr__pnp_05v5_W3p40L3p40
.ends

.subckt XM_bjt sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2]/Emitter
+ VSUBS
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|0] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|1] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|2]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|3] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6|4]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
.ends

.subckt sky130_fd_pr__res_high_po_1p41_GWJZ59 a_n141_n10832# a_n271_n10962# a_n141_10400#
X0 a_n141_n10832# a_n141_10400# a_n271_n10962# sky130_fd_pr__res_high_po_1p41 l=1.04e+08u
.ends

.subckt sky130_fd_pr__res_high_po_1p41_6ZUZ5C a_n271_n1372# a_n141_810# a_n141_n1242#
X0 a_n141_n1242# a_n141_810# a_n271_n1372# sky130_fd_pr__res_high_po_1p41 l=8.1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MUAP4U a_n100_n344# a_n416_118# a_358_118# a_n416_n247#
+ a_n674_118# a_n616_n344# a_n158_118# a_n100_21# a_n358_21# a_158_21# a_358_n247#
+ w_n812_n466# a_158_n344# a_100_n247# a_n674_n247# a_n616_21# a_416_21# a_n158_n247#
+ a_616_118# a_100_118# a_616_n247# a_n358_n344# a_416_n344#
X0 a_100_118# a_n100_21# a_n158_118# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_616_118# a_416_21# a_358_118# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_100_n247# a_n100_n344# a_n158_n247# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_n416_n247# a_n616_n344# a_n674_n247# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_n158_n247# a_n358_n344# a_n416_n247# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X5 a_358_118# a_158_21# a_100_118# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X6 a_n416_118# a_n616_21# a_n674_118# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X7 a_n158_118# a_n358_21# a_n416_118# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X8 a_358_n247# a_158_n344# a_100_n247# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X9 a_616_n247# a_416_n344# a_358_n247# w_n812_n466# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt XM_otabias_pmos m1_143_85# m1_330_160# m1_70_320# sky130_fd_pr__pfet_01v8_lvt_MUAP4U_0/w_n812_n466#
Xsky130_fd_pr__pfet_01v8_lvt_MUAP4U_0 m1_143_85# m1_330_160# m1_70_320# m1_330_160#
+ m1_70_320# m1_143_85# m1_70_320# m1_143_85# m1_143_85# m1_143_85# m1_70_320# sky130_fd_pr__pfet_01v8_lvt_MUAP4U_0/w_n812_n466#
+ m1_143_85# m1_330_160# m1_70_320# m1_143_85# m1_143_85# m1_70_320# m1_330_160# m1_330_160#
+ m1_330_160# m1_143_85# m1_143_85# sky130_fd_pr__pfet_01v8_lvt_MUAP4U
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_9UM225 a_n932_n247# a_n100_n344# a_n416_118# a_674_21#
+ a_n358_386# a_n416_n612# a_874_118# a_358_118# w_n968_18# a_874_n612# a_158_n709#
+ a_n416_n247# w_n968_n712# a_n674_118# w_n968_383# a_n874_n709# a_874_n247# a_416_386#
+ a_n616_n344# a_n158_118# a_n100_21# a_674_n344# w_n968_n347# a_358_n612# a_n358_21#
+ a_100_n612# a_n674_n612# a_158_21# a_n358_n709# a_358_n247# a_616_483# a_100_483#
+ a_674_386# a_158_n344# a_158_386# a_416_n709# a_n100_n709# a_100_n247# a_n674_n247#
+ a_n932_483# a_n616_21# a_n416_483# a_n158_n612# a_n874_n344# a_416_21# a_n100_386#
+ a_n616_386# a_874_483# a_616_n612# a_358_483# a_n158_n247# a_616_118# a_100_118#
+ a_n932_n612# a_n616_n709# a_616_n247# a_n358_n344# a_n674_483# a_674_n709# a_n874_21#
+ a_416_n344# a_n932_118# a_n158_483# a_n874_386#
X0 a_100_118# a_n100_21# a_n158_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X1 a_n158_483# a_n358_386# a_n416_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X2 a_874_483# a_674_386# a_616_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X3 a_874_n247# a_674_n344# a_616_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X4 a_874_n612# a_674_n709# a_616_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X5 a_100_483# a_n100_386# a_n158_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X6 a_n674_118# a_n874_21# a_n932_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X7 a_616_118# a_416_21# a_358_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X8 a_n674_483# a_n874_386# a_n932_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X9 a_100_n247# a_n100_n344# a_n158_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X10 a_100_n612# a_n100_n709# a_n158_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X11 a_n416_n247# a_n616_n344# a_n674_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X12 a_n416_n612# a_n616_n709# a_n674_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X13 a_616_483# a_416_386# a_358_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X14 a_n158_n247# a_n358_n344# a_n416_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X15 a_n158_n612# a_n358_n709# a_n416_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X16 a_358_118# a_158_21# a_100_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X17 a_n416_118# a_n616_21# a_n674_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X18 a_n674_n612# a_n874_n709# a_n932_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X19 a_n674_n247# a_n874_n344# a_n932_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X20 a_358_483# a_158_386# a_100_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X21 a_874_118# a_674_21# a_616_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X22 a_616_n612# a_416_n709# a_358_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=2.9e+11p ps=2.58e+06u w=1e+06u l=1e+06u
X23 a_n416_483# a_n616_386# a_n674_483# w_n968_383# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X24 a_n158_118# a_n358_21# a_n416_118# w_n968_18# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X25 a_358_n247# a_158_n344# a_100_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=0p ps=0u w=1e+06u l=1e+06u
X26 a_616_n247# a_416_n344# a_358_n247# w_n968_n347# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
X27 a_358_n612# a_158_n709# a_100_n612# w_n968_n712# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=1e+06u
.ends

.subckt XM_feedbackmir2 m1_290_100# m1_102_14# m1_102_742# m1_30_240# m1_104_1108#
+ m1_100_382# w_n140_n160#
Xsky130_fd_pr__pfet_01v8_lvt_9UM225_0 m1_30_240# m1_100_382# m1_30_240# m1_102_742#
+ m1_104_1108# m1_30_240# m1_290_100# m1_290_100# w_n140_n160# m1_290_100# m1_102_14#
+ m1_30_240# w_n140_n160# m1_290_100# w_n140_n160# m1_102_14# m1_290_100# m1_104_1108#
+ m1_100_382# m1_290_100# m1_102_742# m1_100_382# w_n140_n160# m1_290_100# m1_102_742#
+ m1_30_240# m1_290_100# m1_102_742# m1_102_14# m1_290_100# m1_30_240# m1_30_240#
+ m1_104_1108# m1_100_382# m1_104_1108# m1_102_14# m1_102_14# m1_30_240# m1_290_100#
+ m1_30_240# m1_102_742# m1_30_240# m1_290_100# m1_100_382# m1_102_742# m1_104_1108#
+ m1_104_1108# m1_290_100# m1_30_240# m1_290_100# m1_290_100# m1_30_240# m1_30_240#
+ m1_30_240# m1_102_14# m1_30_240# m1_100_382# m1_290_100# m1_102_14# m1_102_742#
+ m1_100_382# m1_30_240# m1_290_100# m1_104_1108# sky130_fd_pr__pfet_01v8_lvt_9UM225
.ends

.subckt XM_bjt_out sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2]/Emitter VSUBS
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|0] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|0] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|0] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|1] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|1] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|1] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|2] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2] sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|2]/Emitter
+ VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|2] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|3] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|3] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|3] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0|4] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1|4] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
Xsky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2|4] VSUBS VSUBS VSUBS sky130_fd_pr__rf_pnp_05v5_W3p40L3p40 m=1
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_D74VRS a_n345_118# a_n661_n1247# a_445_118# a_977_n1344#
+ a_n761_1386# a_n819_1483# a_n345_n2612# a_n819_n2612# a_977_21# a_n977_n1247# a_n345_1483#
+ a_187_21# a_n187_118# a_287_118# a_n187_n2612# a_n1135_1483# a_n977_1483# a_n661_n2612#
+ a_n445_21# a_n819_118# a_n503_1483# a_129_1483# a_919_118# a_n977_n2612# a_n1077_21#
+ a_n661_118# a_761_118# a_29_21# a_345_21# a_29_n2709# a_n661_1483# a_287_1483# a_n603_21#
+ a_29_n1344# a_129_n1247# a_29_1386# a_919_1483# a_603_n1247# a_n129_1386# a_445_1483#
+ a_187_1386# a_n1135_118# a_445_n1247# a_n129_n2709# w_n1273_n2831# a_503_21# a_919_n1247#
+ a_1077_n1247# a_129_n2612# a_1077_1483# a_n603_n2709# a_287_n1247# a_n287_1386#
+ a_n129_n1344# a_819_1386# a_n1077_n2709# a_n977_118# a_1077_118# a_603_n2612# a_n1077_1386#
+ a_603_1483# a_761_n1247# a_n445_n2709# a_503_n2709# a_n29_n1247# a_n919_21# a_n919_n2709#
+ a_345_1386# a_n603_n1344# a_n761_21# a_n129_21# a_129_118# a_445_n2612# a_n919_1386#
+ a_n1077_n1344# a_n287_n2709# a_345_n2709# a_919_n2612# a_819_n2709# a_503_n1344#
+ a_1077_n2612# a_977_1386# a_n445_n1344# a_n445_1386# a_n919_n1344# a_761_1483# a_n1135_n1247#
+ a_n761_n2709# a_287_n2612# a_187_n2709# a_819_21# a_n503_n1247# a_661_21# a_345_n1344#
+ a_n29_118# a_n287_n1344# a_819_n1344# a_503_1386# a_761_n2612# a_n29_1483# a_661_n2709#
+ a_n29_n2612# a_n503_118# a_n761_n1344# a_n345_n1247# a_603_118# a_187_n1344# a_n819_n1247#
+ a_n603_1386# a_n187_1483# a_977_n2709# a_661_n1344# a_n187_n1247# a_661_1386# a_n1135_n2612#
+ a_n287_21# a_n503_n2612#
X0 a_n819_n1247# a_n919_n1344# a_n977_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X1 a_n977_n1247# a_n1077_n1344# a_n1135_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X2 a_603_n2612# a_503_n2709# a_445_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X3 a_n977_118# a_n1077_21# a_n1135_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X4 a_603_n1247# a_503_n1344# a_445_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X5 a_761_n2612# a_661_n2709# a_603_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X6 a_n819_1483# a_n919_1386# a_n977_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X7 a_761_n1247# a_661_n1344# a_603_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X8 a_n661_1483# a_n761_1386# a_n819_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X9 a_919_1483# a_819_1386# a_761_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X10 a_n187_1483# a_n287_1386# a_n345_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X11 a_761_1483# a_661_1386# a_603_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X12 a_n661_118# a_n761_21# a_n819_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X13 a_n503_n2612# a_n603_n2709# a_n661_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X14 a_129_118# a_29_21# a_n29_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X15 a_287_n2612# a_187_n2709# a_129_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X16 a_n187_118# a_n287_21# a_n345_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X17 a_n503_n1247# a_n603_n1344# a_n661_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X18 a_n661_n2612# a_n761_n2709# a_n819_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X19 a_287_1483# a_187_1386# a_129_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X20 a_n661_n1247# a_n761_n1344# a_n819_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X21 a_287_n1247# a_187_n1344# a_129_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X22 a_n819_118# a_n919_21# a_n977_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X23 a_n345_118# a_n445_21# a_n503_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X24 a_n503_118# a_n603_21# a_n661_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X25 a_n29_n2612# a_n129_n2709# a_n187_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X26 a_n345_1483# a_n445_1386# a_n503_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X27 a_n29_n1247# a_n129_n1344# a_n187_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X28 a_n187_n2612# a_n287_n2709# a_n345_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X29 a_n29_118# a_n129_21# a_n187_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X30 a_129_1483# a_29_1386# a_n29_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X31 a_n187_n1247# a_n287_n1344# a_n345_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X32 a_445_1483# a_345_1386# a_287_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X33 a_1077_118# a_977_21# a_919_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X34 a_129_n2612# a_29_n2709# a_n29_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X35 a_n977_1483# a_n1077_1386# a_n1135_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X36 a_129_n1247# a_29_n1344# a_n29_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X37 a_445_n2612# a_345_n2709# a_287_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X38 a_n503_1483# a_n603_1386# a_n661_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X39 a_1077_1483# a_977_1386# a_919_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X40 a_761_118# a_661_21# a_603_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X41 a_287_118# a_187_21# a_129_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X42 a_445_n1247# a_345_n1344# a_287_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X43 a_919_n2612# a_819_n2709# a_761_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X44 a_n29_1483# a_n129_1386# a_n187_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X45 a_603_1483# a_503_1386# a_445_1483# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X46 a_445_118# a_345_21# a_287_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X47 a_919_118# a_819_21# a_761_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X48 a_919_n1247# a_819_n1344# a_761_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X49 a_1077_n2612# a_977_n2709# a_919_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X50 a_1077_n1247# a_977_n1344# a_919_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=1.74e+12p pd=1.258e+07u as=0p ps=0u w=6e+06u l=500000u
X51 a_603_118# a_503_21# a_445_118# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X52 a_n345_n2612# a_n445_n2709# a_n503_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X53 a_n345_n1247# a_n445_n1344# a_n503_n1247# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=6e+06u l=500000u
X54 a_n819_n2612# a_n919_n2709# a_n977_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
X55 a_n977_n2612# a_n1077_n2709# a_n1135_n2612# w_n1273_n2831# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=1.74e+12p ps=1.258e+07u w=6e+06u l=500000u
.ends

.subckt XM_cs li_876_5462# m1_52_164# m1_147_79#
Xsky130_fd_pr__pfet_01v8_lvt_D74VRS_0 li_876_5462# li_876_5462# m1_52_164# m1_147_79#
+ m1_147_79# m1_52_164# li_876_5462# m1_52_164# m1_147_79# li_876_5462# li_876_5462#
+ m1_147_79# m1_52_164# li_876_5462# m1_52_164# m1_52_164# li_876_5462# li_876_5462#
+ m1_147_79# m1_52_164# m1_52_164# m1_52_164# li_876_5462# li_876_5462# m1_147_79#
+ li_876_5462# m1_52_164# m1_147_79# m1_147_79# m1_147_79# li_876_5462# li_876_5462#
+ m1_147_79# m1_147_79# m1_52_164# m1_147_79# li_876_5462# li_876_5462# m1_147_79#
+ m1_52_164# m1_147_79# m1_52_164# m1_52_164# m1_147_79# li_876_5462# m1_147_79# li_876_5462#
+ m1_52_164# m1_52_164# m1_52_164# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_147_79#
+ m1_147_79# li_876_5462# m1_52_164# li_876_5462# m1_147_79# li_876_5462# m1_52_164#
+ m1_147_79# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_147_79# m1_147_79# m1_147_79#
+ m1_147_79# m1_52_164# m1_52_164# m1_147_79# m1_147_79# m1_147_79# m1_147_79# li_876_5462#
+ m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_147_79# m1_147_79# m1_147_79# m1_52_164#
+ m1_52_164# m1_147_79# li_876_5462# m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_147_79#
+ li_876_5462# m1_147_79# m1_147_79# m1_147_79# m1_52_164# li_876_5462# m1_147_79#
+ li_876_5462# m1_52_164# m1_147_79# li_876_5462# li_876_5462# m1_147_79# m1_52_164#
+ m1_147_79# m1_52_164# m1_147_79# m1_147_79# m1_52_164# m1_147_79# m1_52_164# m1_147_79#
+ m1_52_164# sky130_fd_pr__pfet_01v8_lvt_D74VRS
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_E96B6C a_29_n507# a_n287_n419# a_n229_n507# a_287_n507#
+ a_229_n419# a_n545_n419# a_n487_n507# a_n29_n419# a_487_n419# VSUBS
X0 a_487_n419# a_287_n507# a_229_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X1 a_n29_n419# a_n229_n507# a_n287_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X2 a_229_n419# a_29_n507# a_n29_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=4.5e+06u l=1e+06u
X3 a_n287_n419# a_n487_n507# a_n545_n419# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_A5VCMN a_229_n481# a_29_n507# a_n545_n481# a_n229_n507#
+ a_287_n507# a_n29_n481# a_487_n481# a_n487_n507# a_n287_n481# VSUBS
X0 a_487_n481# a_287_n507# a_229_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=1.305e+12p pd=9.58e+06u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X1 a_229_n481# a_29_n507# a_n29_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X2 a_n29_n481# a_n229_n507# a_n287_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
X3 a_n287_n481# a_n487_n507# a_n545_n481# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=1.305e+12p ps=9.58e+06u w=4.5e+06u l=1e+06u
.ends

.subckt XM_diffpair m1_160_200# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS m1_30_1280#
+ m1_30_n1060# m1_280_n670# m1_551_360#
Xsky130_fd_pr__nfet_01v8_lvt_E96B6C_0 m1_551_360# m1_280_n670# m1_551_360# m1_160_200#
+ m1_280_n670# m1_30_1280# m1_160_200# m1_30_n1060# m1_30_1280# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_E96B6C
Xsky130_fd_pr__nfet_01v8_lvt_A5VCMN_0 m1_280_n670# m1_160_200# m1_30_n1060# m1_160_200#
+ m1_551_360# m1_30_1280# m1_30_n1060# m1_551_360# m1_280_n670# sky130_fd_pr__nfet_01v8_lvt_E96B6C_0/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_A5VCMN
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_EN3Q86 c1_n1650_n2140# m3_n1750_n2240#
X0 c1_n1650_n2140# m3_n1750_n2240# sky130_fd_pr__cap_mim_m3_1 l=2.14e+07u w=1.6e+07u
.ends

.subckt sky130_fd_pr__res_high_po_2p85_7J2RPB a_n285_n1642# a_n415_n1772# a_n285_1210#
X0 a_n285_n1642# a_n285_1210# a_n415_n1772# sky130_fd_pr__res_high_po_2p85 l=1.21e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_USQY94 a_n1174_n1403# a_658_109# a_n716_n1403#
+ a_200_109# a_n1116_21# a_1116_865# a_n258_n1403# a_n200_n1491# a_716_n1491# a_n1174_n647#
+ a_n200_21# a_n658_n1491# a_n200_n735# a_n258_865# a_1116_109# a_200_n647# a_258_21#
+ a_n658_21# a_1116_n1403# a_258_n1491# a_258_777# a_n1276_n1577# a_n1116_n735# a_n258_109#
+ a_n716_n647# a_n1174_865# a_n658_777# a_n200_777# a_n258_n647# a_n716_865# a_n658_n735#
+ a_200_n1403# a_1116_n647# a_n1174_109# a_716_21# a_658_n1403# a_716_n735# a_658_865#
+ a_716_777# a_658_n647# a_258_n735# a_200_865# a_n1116_n1491# a_n716_109# a_n1116_777#
X0 a_658_n1403# a_258_n1491# a_200_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X1 a_n716_n1403# a_n1116_n1491# a_n1174_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X2 a_658_109# a_258_21# a_200_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X3 a_1116_n647# a_716_n735# a_658_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X4 a_1116_n1403# a_716_n1491# a_658_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X5 a_200_865# a_n200_777# a_n258_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X6 a_1116_109# a_716_21# a_658_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X7 a_200_n647# a_n200_n735# a_n258_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X8 a_n716_n647# a_n1116_n735# a_n1174_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X9 a_n258_865# a_n658_777# a_n716_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X10 a_n716_865# a_n1116_777# a_n1174_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X11 a_658_n647# a_258_n735# a_200_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X12 a_200_109# a_n200_21# a_n258_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X13 a_658_865# a_258_777# a_200_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X14 a_n258_109# a_n658_21# a_n716_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X15 a_n258_n647# a_n658_n735# a_n716_n647# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
X16 a_200_n1403# a_n200_n1491# a_n258_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X17 a_1116_865# a_716_777# a_658_865# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=8.7e+11p pd=6.58e+06u as=0p ps=0u w=3e+06u l=2e+06u
X18 a_n716_109# a_n1116_21# a_n1174_109# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=8.7e+11p ps=6.58e+06u w=3e+06u l=2e+06u
X19 a_n258_n1403# a_n658_n1491# a_n716_n1403# a_n1276_n1577# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3e+06u l=2e+06u
.ends

.subckt XM_actload2 m1_985_79# m1_522_658# m1_522_1414# m1_62_1668# m1_522_2926# m1_520_2170#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_USQY94_0 m1_62_1668# m1_62_1668# m1_522_658# m1_520_2170#
+ m1_985_79# m1_522_2926# m1_62_1668# m1_985_79# m1_985_79# m1_62_1668# m1_985_79#
+ m1_985_79# m1_985_79# m1_62_1668# m1_520_2170# m1_522_1414# m1_985_79# m1_985_79#
+ m1_522_658# m1_985_79# m1_985_79# VSUBS m1_985_79# m1_62_1668# m1_522_1414# m1_62_1668#
+ m1_985_79# m1_985_79# m1_62_1668# m1_522_2926# m1_985_79# m1_522_658# m1_522_1414#
+ m1_62_1668# m1_985_79# m1_62_1668# m1_985_79# m1_62_1668# m1_985_79# m1_62_1668#
+ m1_985_79# m1_522_2926# m1_985_79# m1_520_2170# m1_985_79# sky130_fd_pr__nfet_01v8_lvt_USQY94
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_7MFZYU a_n429_299# a_29_299# a_n487_n725# a_429_387#
+ a_429_n1281# a_n29_n725# a_n487_943# a_n429_n813# a_429_n725# a_n487_n169# a_29_n813#
+ a_n29_943# a_n589_n1455# a_29_n1369# a_n29_n1281# a_n29_n169# a_n487_387# a_n429_n257#
+ a_29_855# a_n429_855# a_n429_n1369# a_429_n169# a_n487_n1281# a_29_n257# a_n29_387#
+ a_429_943#
X0 a_429_n169# a_29_n257# a_n29_n169# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X1 a_429_n725# a_29_n813# a_n29_n725# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X2 a_n29_n1281# a_n429_n1369# a_n487_n1281# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X3 a_429_387# a_29_299# a_n29_387# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X4 a_429_943# a_29_855# a_n29_943# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X5 a_429_n1281# a_29_n1369# a_n29_n1281# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=2e+06u
X6 a_n29_n169# a_n429_n257# a_n487_n169# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X7 a_n29_n725# a_n429_n813# a_n487_n725# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X8 a_n29_943# a_n429_855# a_n487_943# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
X9 a_n29_387# a_n429_299# a_n487_387# a_n589_n1455# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=2e+06u
.ends

.subckt XM_tail m1_530_330# m1_780_80# VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_7MFZYU_0 m1_780_80# m1_780_80# VSUBS VSUBS VSUBS m1_530_330#
+ VSUBS m1_780_80# VSUBS VSUBS m1_780_80# m1_530_330# VSUBS m1_780_80# m1_530_330#
+ m1_530_330# VSUBS m1_780_80# m1_780_80# m1_780_80# m1_780_80# VSUBS VSUBS m1_780_80#
+ m1_530_330# VSUBS sky130_fd_pr__nfet_01v8_lvt_7MFZYU
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_MBDTEX a_745_n236# a_545_n262# a_1777_n236# a_1577_n262#
+ a_229_n236# a_n1577_n236# a_2035_n236# a_n1777_n262# a_29_n262# w_n2129_n298# a_n545_n236#
+ a_n745_n262# a_1003_n236# a_803_n262# a_n2035_n262# a_1835_n262# a_n29_n236# a_n229_n262#
+ a_487_n236# a_287_n262# a_n1003_n262# a_n1835_n236# a_n803_n236# a_1519_n236# a_n2093_n236#
+ a_1319_n262# a_1261_n236# a_1061_n262# a_n1319_n236# a_n287_n236# a_n1061_n236#
+ a_n1519_n262# a_n487_n262# a_n1261_n262#
X0 a_n1061_n236# a_n1261_n262# a_n1319_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_745_n236# a_545_n262# a_487_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X2 a_1003_n236# a_803_n262# a_745_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X3 a_487_n236# a_287_n262# a_229_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X4 a_2035_n236# a_1835_n262# a_1777_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X5 a_1777_n236# a_1577_n262# a_1519_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X6 a_1261_n236# a_1061_n262# a_1003_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X7 a_n1835_n236# a_n2035_n262# a_n2093_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X8 a_n29_n236# a_n229_n262# a_n287_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X9 a_229_n236# a_29_n262# a_n29_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X10 a_n1319_n236# a_n1519_n262# a_n1577_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X11 a_n545_n236# a_n745_n262# a_n803_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X12 a_n803_n236# a_n1003_n262# a_n1061_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X13 a_n287_n236# a_n487_n262# a_n545_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_n1577_n236# a_n1777_n262# a_n1835_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 a_1519_n236# a_1319_n262# a_1261_n236# w_n2129_n298# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_B64SAM a_545_n261# a_1777_n164# a_1577_n261# a_229_n164#
+ a_n1577_n164# a_2035_n164# a_n545_n164# a_29_n261# a_n1777_n261# a_n745_n261# a_1003_n164#
+ a_803_n261# a_n2035_n261# a_n29_n164# a_487_n164# a_1835_n261# a_n229_n261# w_n2129_n264#
+ a_n1835_n164# a_287_n261# a_n1003_n261# a_n803_n164# a_1519_n164# a_n2093_n164#
+ a_1261_n164# a_1319_n261# a_n1319_n164# a_1061_n261# a_n287_n164# a_n1061_n164#
+ a_n1519_n261# a_745_n164# a_n487_n261# a_n1261_n261#
X0 a_n29_n164# a_n229_n261# a_n287_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X1 a_229_n164# a_29_n261# a_n29_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X2 a_n1319_n164# a_n1519_n261# a_n1577_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X3 a_n545_n164# a_n745_n261# a_n803_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X4 a_n287_n164# a_n487_n261# a_n545_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X5 a_n803_n164# a_n1003_n261# a_n1061_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X6 a_n1577_n164# a_n1777_n261# a_n1835_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X7 a_1519_n164# a_1319_n261# a_1261_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X8 a_n1061_n164# a_n1261_n261# a_n1319_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X9 a_1003_n164# a_803_n261# a_745_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X10 a_745_n164# a_545_n261# a_487_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
X11 a_487_n164# a_287_n261# a_229_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X12 a_1777_n164# a_1577_n261# a_1519_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X13 a_2035_n164# a_1835_n261# a_1777_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=5.8e+11p pd=4.58e+06u as=0p ps=0u w=2e+06u l=1e+06u
X14 a_1261_n164# a_1061_n261# a_1003_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=2e+06u l=1e+06u
X15 a_n1835_n164# a_n2035_n261# a_n2093_n164# w_n2129_n264# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=5.8e+11p ps=4.58e+06u w=2e+06u l=1e+06u
.ends

.subckt XM_ppair w_n220_n1060# m1_240_n480# m1_70_n360#
Xsky130_fd_pr__pfet_01v8_lvt_MBDTEX_0 m1_70_n360# m1_70_n360# m1_240_n480# m1_70_n360#
+ m1_240_n480# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# w_n220_n1060# w_n220_n1060#
+ m1_70_n360# w_n220_n1060# m1_70_n360# m1_70_n360# m1_70_n360# w_n220_n1060# m1_70_n360#
+ w_n220_n1060# m1_70_n360# m1_70_n360# m1_240_n480# m1_70_n360# w_n220_n1060# w_n220_n1060#
+ m1_70_n360# m1_70_n360# m1_70_n360# m1_70_n360# m1_240_n480# w_n220_n1060# m1_70_n360#
+ m1_70_n360# m1_70_n360# sky130_fd_pr__pfet_01v8_lvt_MBDTEX
Xsky130_fd_pr__pfet_01v8_lvt_B64SAM_0 m1_70_n360# m1_70_n360# m1_70_n360# m1_70_n360#
+ w_n220_n1060# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# m1_70_n360# w_n220_n1060#
+ m1_70_n360# m1_70_n360# w_n220_n1060# w_n220_n1060# m1_70_n360# m1_70_n360# w_n220_n1060#
+ m1_70_n360# m1_70_n360# m1_70_n360# m1_240_n480# w_n220_n1060# w_n220_n1060# m1_240_n480#
+ m1_70_n360# m1_240_n480# m1_70_n360# m1_70_n360# w_n220_n1060# m1_70_n360# m1_240_n480#
+ m1_70_n360# m1_70_n360# sky130_fd_pr__pfet_01v8_lvt_B64SAM
.ends

.subckt opamp_realcomp3_usefinger in_n in_p out bias_0p7 vdd vss
XXM_cs_0 vdd out first_stage_out XM_cs
XXM_diffpair_0 in_p vss first_stage_out ppair_gate m2_n4080_2260# in_n XM_diffpair
Xsky130_fd_pr__cap_mim_m3_1_EN3Q86_0 first_stage_out m1_6290_1100# sky130_fd_pr__cap_mim_m3_1_EN3Q86
Xsky130_fd_pr__res_high_po_2p85_7J2RPB_0 out vss m1_6290_1100# sky130_fd_pr__res_high_po_2p85_7J2RPB
XXM_actload2_0 bias_0p7 out out vss out out vss XM_actload2
XXM_tail_0 m2_n4080_2260# bias_0p7 vss XM_tail
XXM_ppair_0 vdd first_stage_out ppair_gate XM_ppair
.ends

.subckt sky130_fd_pr__res_high_po_1p41_HX7ZEK a_n271_n5312# a_n141_n5182# a_n141_4750#
X0 a_n141_n5182# a_n141_4750# a_n271_n5312# sky130_fd_pr__res_high_po_1p41 l=4.75e+07u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_QA4PPD li_n560_n643# a_n458_n469# a_n400_n557#
+ a_400_n469# a_n560_n643#
X0 a_400_n469# a_n400_n557# a_n458_n469# a_n560_n643# sky130_fd_pr__nfet_01v8_lvt ad=1.45e+12p pd=1.058e+07u as=1.45e+12p ps=1.058e+07u w=5e+06u l=4e+06u
.ends

.subckt XM_otabias_nmos sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_n458_n469# sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/li_n560_n643#
+ sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_n400_n557# sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_400_n469#
+ VSUBS
Xsky130_fd_pr__nfet_01v8_lvt_QA4PPD_0 sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/li_n560_n643#
+ sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_n458_n469# sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_n400_n557#
+ sky130_fd_pr__nfet_01v8_lvt_QA4PPD_0/a_400_n469# VSUBS sky130_fd_pr__nfet_01v8_lvt_QA4PPD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_64DJ5N a_n945_n831# a_n487_n831# a_n29_n831# a_887_n831#
+ a_n887_n857# a_429_n831# a_n429_n857# a_487_n857# a_29_n857# VSUBS
X0 a_429_n831# a_29_n857# a_n29_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X1 a_887_n831# a_487_n857# a_429_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=2e+06u
X2 a_n487_n831# a_n887_n857# a_n945_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X3 a_n29_n831# a_n429_n857# a_n487_n831# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_64S6GM a_n945_n769# a_n487_n769# a_n887_n857#
+ a_n29_n769# a_887_n769# a_n429_n857# a_487_n857# a_429_n769# a_29_n857# VSUBS
X0 a_429_n769# a_29_n857# a_n29_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X1 a_887_n769# a_487_n857# a_429_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=0p ps=0u w=8e+06u l=2e+06u
X2 a_n487_n769# a_n887_n857# a_n945_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=2.32e+12p pd=1.658e+07u as=2.32e+12p ps=1.658e+07u w=8e+06u l=2e+06u
X3 a_n29_n769# a_n429_n857# a_n487_n769# VSUBS sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=8e+06u l=2e+06u
.ends

.subckt XM_output_mirr sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS m1_62_n98# m1_62_n3610#
+ m1_n10_n960# m1_n10_n4460# m1_450_n4460#
Xsky130_fd_pr__nfet_01v8_lvt_64DJ5N_0 m1_n10_n960# m1_450_n4460# m1_n10_n960# m1_n10_n960#
+ m1_62_n98# m1_450_n4460# m1_62_n98# m1_62_n98# m1_62_n98# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64DJ5N
Xsky130_fd_pr__nfet_01v8_lvt_64DJ5N_1 m1_n10_n4460# m1_450_n4460# m1_n10_n4460# m1_n10_n4460#
+ m1_62_n3610# m1_450_n4460# m1_62_n3610# m1_62_n3610# m1_62_n3610# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64DJ5N
Xsky130_fd_pr__nfet_01v8_lvt_64S6GM_0 m1_n10_n960# m1_450_n4460# m1_62_n98# m1_n10_n960#
+ m1_n10_n960# m1_62_n98# m1_62_n98# m1_450_n4460# m1_62_n98# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64S6GM
Xsky130_fd_pr__nfet_01v8_lvt_64S6GM_1 m1_n10_n4460# m1_450_n4460# m1_62_n3610# m1_n10_n4460#
+ m1_n10_n4460# m1_62_n3610# m1_62_n3610# m1_450_n4460# m1_62_n3610# sky130_fd_pr__nfet_01v8_lvt_64S6GM_1/VSUBS
+ sky130_fd_pr__nfet_01v8_lvt_64S6GM
.ends

.subckt XM_output_mirr_combined XM_output_mirr_7/m1_450_n4460# XM_output_mirr_7/m1_62_n98#
+ XM_output_mirr_2/m1_n10_n4460# XM_output_mirr_2/m1_62_n98# XM_output_mirr_2/m1_n10_n960#
+ XM_output_mirr_4/m1_n10_n960# XM_output_mirr_7/m1_62_n3610# XM_output_mirr_2/m1_450_n4460#
+ XM_output_mirr_4/m1_62_n98# XM_output_mirr_2/m1_62_n3610# XM_output_mirr_0/m1_450_n4460#
+ XM_output_mirr_5/m1_62_n98# XM_output_mirr_0/m1_62_n98# XM_output_mirr_6/m1_62_n3610#
+ XM_output_mirr_5/m1_n10_n4460# XM_output_mirr_3/m1_n10_n4460# XM_output_mirr_5/m1_62_n3610#
+ XM_output_mirr_6/m1_450_n4460# XM_output_mirr_3/m1_450_n4460# XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr_7/m1_n10_n960# XM_output_mirr_0/m1_62_n3610# XM_output_mirr_3/m1_62_n98#
+ XM_output_mirr_6/m1_n10_n4460# XM_output_mirr_5/m1_450_n4460# XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr_1/m1_n10_n960# XM_output_mirr_6/m1_62_n98# XM_output_mirr_3/m1_62_n3610#
+ XM_output_mirr_6/m1_n10_n960# XM_output_mirr_5/m1_n10_n960# XM_output_mirr_7/m1_n10_n4460#
+ XM_output_mirr_1/m1_n10_n4460# XM_output_mirr_1/m1_62_n98# XM_output_mirr_4/m1_62_n3610#
+ XM_output_mirr_4/m1_n10_n4460# XM_output_mirr_0/m1_n10_n960# XM_output_mirr_0/m1_n10_n4460#
+ XM_output_mirr_1/m1_62_n3610# VSUBS XM_output_mirr_3/m1_n10_n960#
XXM_output_mirr_0 VSUBS XM_output_mirr_0/m1_62_n98# XM_output_mirr_0/m1_62_n3610#
+ XM_output_mirr_0/m1_n10_n960# XM_output_mirr_0/m1_n10_n4460# XM_output_mirr_0/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_1 VSUBS XM_output_mirr_1/m1_62_n98# XM_output_mirr_1/m1_62_n3610#
+ XM_output_mirr_1/m1_n10_n960# XM_output_mirr_1/m1_n10_n4460# XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_2 VSUBS XM_output_mirr_2/m1_62_n98# XM_output_mirr_2/m1_62_n3610#
+ XM_output_mirr_2/m1_n10_n960# XM_output_mirr_2/m1_n10_n4460# XM_output_mirr_2/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_3 VSUBS XM_output_mirr_3/m1_62_n98# XM_output_mirr_3/m1_62_n3610#
+ XM_output_mirr_3/m1_n10_n960# XM_output_mirr_3/m1_n10_n4460# XM_output_mirr_3/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_4 VSUBS XM_output_mirr_4/m1_62_n98# XM_output_mirr_4/m1_62_n3610#
+ XM_output_mirr_4/m1_n10_n960# XM_output_mirr_4/m1_n10_n4460# XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_5 VSUBS XM_output_mirr_5/m1_62_n98# XM_output_mirr_5/m1_62_n3610#
+ XM_output_mirr_5/m1_n10_n960# XM_output_mirr_5/m1_n10_n4460# XM_output_mirr_5/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_6 VSUBS XM_output_mirr_6/m1_62_n98# XM_output_mirr_6/m1_62_n3610#
+ XM_output_mirr_6/m1_n10_n960# XM_output_mirr_6/m1_n10_n4460# XM_output_mirr_6/m1_450_n4460#
+ XM_output_mirr
XXM_output_mirr_7 VSUBS XM_output_mirr_7/m1_62_n98# XM_output_mirr_7/m1_62_n3610#
+ XM_output_mirr_7/m1_n10_n960# XM_output_mirr_7/m1_n10_n4460# XM_output_mirr_7/m1_450_n4460#
+ XM_output_mirr
.ends

.subckt XM_output_mirr_combined_with_dummy XM_output_mirr_combined_0/XM_output_mirr_5/m1_n10_n960#
+ m1_300_5420# XM_output_mirr_combined_0/XM_output_mirr_4/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_3/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_7/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_2/m1_n10_n960#
+ m2_300_360# XM_output_mirr_combined_0/XM_output_mirr_6/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_1/m1_n10_n960#
+ VSUBS
XXM_output_mirr_combined_0 XM_output_mirr_combined_0/XM_output_mirr_7/m1_450_n4460#
+ m1_300_5420# m2_300_360# m1_300_5420# XM_output_mirr_combined_0/XM_output_mirr_2/m1_n10_n960#
+ XM_output_mirr_combined_0/XM_output_mirr_4/m1_n10_n960# m1_740_1920# XM_output_mirr_combined_0/XM_output_mirr_2/m1_450_n4460#
+ m1_300_5420# m1_740_1920# m1_740_1920# m1_300_5420# m1_300_5420# m1_740_1920# m2_300_360#
+ m2_300_360# m1_740_1920# XM_output_mirr_combined_0/XM_output_mirr_6/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_3/m1_450_n4460# XM_output_mirr_combined_0/XM_output_mirr_4/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_7/m1_n10_n960# m1_740_1920# m1_300_5420#
+ m2_300_360# XM_output_mirr_combined_0/XM_output_mirr_5/m1_450_n4460# XM_output_mirr_combined_0/XM_output_mirr_1/m1_450_n4460#
+ XM_output_mirr_combined_0/XM_output_mirr_1/m1_n10_n960# m1_300_5420# m1_740_1920#
+ XM_output_mirr_combined_0/XM_output_mirr_6/m1_n10_n960# XM_output_mirr_combined_0/XM_output_mirr_5/m1_n10_n960#
+ m2_300_360# m2_300_360# m1_300_5420# m1_740_1920# m2_300_360# m1_300_5420# m2_300_360#
+ m1_740_1920# VSUBS XM_output_mirr_combined_0/XM_output_mirr_3/m1_n10_n960# XM_output_mirr_combined
XXM_output_mirr_combined_1 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_2 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_3 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_4 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_5 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_6 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_7 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
XXM_output_mirr_combined_8 VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS VSUBS
+ VSUBS VSUBS VSUBS XM_output_mirr_combined
.ends

.subckt BGR_lvs Iout0 Iout1 Iout2 porst vbg Iout3 Iout4 Iout5 Iout6 VDD VSS
XXM_Rref_0 VSS vd4 VSS XM_Rref
Xsky130_fd_pr__res_high_po_1p41_S8KB58_0 vbg vbe3 VSS sky130_fd_pr__res_high_po_1p41_S8KB58
XXM_pdn_0 VSS vgate porst VDD VSS VSS XM_pdn
XXM_current_gate_with_dummy_0 VDD VDD VDD VDD opamp_realcomp3_usefinger_1/out VDD
+ VDD voutb2 VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD VDD vd4 VDD VDD
+ VDD VDD XM_current_gate_with_dummy
XXM_feedbackmir_0 VDD VDD opamp_realcomp3_usefinger_0/in_n vb vgate XM_feedbackmir
XXM_bjt_0 vbneg opamp_realcomp3_usefinger_0/in_n VSS XM_bjt
Xsky130_fd_pr__res_high_po_1p41_GWJZ59_0 VSS VSS m1_n1770_n3060# sky130_fd_pr__res_high_po_1p41_GWJZ59
Xsky130_fd_pr__res_high_po_1p41_6ZUZ5C_0 VSS vbneg vb sky130_fd_pr__res_high_po_1p41_6ZUZ5C
XXM_otabias_pmos_0 vgate Vota_bias1 VDD VDD XM_otabias_pmos
XXM_feedbackmir2_0 vbg vgate vgate VDD vgate vgate VDD XM_feedbackmir2
XXM_bjt_out_0 vbe3 VSS XM_bjt_out
Xopamp_realcomp3_usefinger_0 opamp_realcomp3_usefinger_0/in_n vb vgate Vota_bias1
+ VDD VSS opamp_realcomp3_usefinger
Xopamp_realcomp3_usefinger_1 vbg vd4 opamp_realcomp3_usefinger_1/out Vota_bias1 VDD
+ VSS opamp_realcomp3_usefinger
Xsky130_fd_pr__res_high_po_1p41_HX7ZEK_0 VSS m1_n1770_n3060# vd4 sky130_fd_pr__res_high_po_1p41_HX7ZEK
XXM_otabias_nmos_0 Vota_bias1 VSS Vota_bias1 VSS VSS XM_otabias_nmos
XXM_output_mirr_combined_with_dummy_0 Iout4 voutb2 Iout3 Iout2 Iout6 Iout1 VSS Iout5
+ Iout0 VSS XM_output_mirr_combined_with_dummy
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_FKGFGD a_1791_122# a_447_122# a_n1905_n100# a_n2433_122#
+ a_591_n100# a_n657_n100# a_n225_n188# a_1407_122# a_2271_n188# a_n321_122# a_207_n100#
+ a_1743_n100# a_927_n188# a_1359_n100# a_2703_n100# a_1311_n188# a_2751_122# a_2319_n100#
+ a_n2577_n100# a_n1185_n188# a_n1665_122# a_n2145_n188# a_n1617_n100# a_n3059_n274#
+ a_n753_n100# a_n369_n100# a_303_n100# a_1455_n100# a_2415_n100# a_639_122# a_1983_122#
+ a_n2673_n100# a_n2289_n100# a_n2625_122# a_n1713_n100# a_n1329_n100# a_n465_n100#
+ a_n897_122# a_n513_122# a_1551_n100# a_n33_n188# a_735_n188# a_1167_n100# a_2511_n100#
+ a_1887_n188# a_2127_n100# a_2847_n188# a_n2385_n100# a_n1857_122# a_15_n100# a_n1425_n100#
+ a_n561_n100# a_831_122# a_n177_n100# a_111_n100# a_879_n100# a_1263_n100# a_2223_n100#
+ a_n2481_n100# a_n2817_122# a_n2097_n100# a_2175_122# a_n2957_n100# a_n1521_n100#
+ a_n1137_n100# a_n1089_122# a_n273_n100# a_n705_122# a_n993_n188# a_975_n100# a_543_n188#
+ a_1695_n188# a_n609_n188# a_159_n188# a_2655_n188# a_n2193_n100# a_1023_122# a_n1233_n100#
+ a_n2049_122# a_n1953_n188# a_n1569_n188# a_n2913_n188# a_63_122# a_n2529_n188# a_687_n100#
+ a_n1281_122# a_1071_n100# a_2031_n100# a_2799_n100# a_2367_122# a_1839_n100# a_255_122#
+ a_n81_n100# a_783_n100# a_n2241_122# a_n849_n100# a_399_n100# a_n801_n188# a_351_n188#
+ a_n417_n188# a_2895_n100# a_1599_122# a_2463_n188# a_1215_122# a_2079_n188# a_1935_n100#
+ a_1503_n188# a_n1041_n100# a_1119_n188# a_n2001_n100# a_n1761_n188# a_n2769_n100#
+ a_n1377_n188# a_n2721_n188# a_n2337_n188# a_n129_122# a_n1809_n100# a_n1473_122#
+ a_n945_n100# a_495_n100# a_2559_122# a_1647_n100# a_2607_n100# a_n2865_n100#
X0 a_n2481_n100# a_n2529_n188# a_n2577_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_n2385_n100# a_n2433_122# a_n2481_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X2 a_n2193_n100# a_n2241_122# a_n2289_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n2097_n100# a_n2145_n188# a_n2193_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X4 a_n2001_n100# a_n2049_122# a_n2097_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_n2673_n100# a_n2721_n188# a_n2769_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_n2577_n100# a_n2625_122# a_n2673_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X7 a_n2289_n100# a_n2337_n188# a_n2385_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X8 a_2031_n100# a_1983_122# a_1935_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X9 a_207_n100# a_159_n188# a_111_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X10 a_303_n100# a_255_122# a_207_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_399_n100# a_351_n188# a_303_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X12 a_495_n100# a_447_122# a_399_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X13 a_591_n100# a_543_n188# a_495_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X14 a_687_n100# a_639_122# a_591_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X15 a_783_n100# a_735_n188# a_687_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X16 a_879_n100# a_831_122# a_783_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X17 a_975_n100# a_927_n188# a_879_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X18 a_n1521_n100# a_n1569_n188# a_n1617_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X19 a_n1425_n100# a_n1473_122# a_n1521_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X20 a_n1233_n100# a_n1281_122# a_n1329_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X21 a_n1137_n100# a_n1185_n188# a_n1233_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X22 a_n1041_n100# a_n1089_122# a_n1137_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X23 a_n1905_n100# a_n1953_n188# a_n2001_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X24 a_n1809_n100# a_n1857_122# a_n1905_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X25 a_n1713_n100# a_n1761_n188# a_n1809_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_n1617_n100# a_n1665_122# a_n1713_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_n1329_n100# a_n1377_n188# a_n1425_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X28 a_n561_n100# a_n609_n188# a_n657_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X29 a_1071_n100# a_1023_122# a_975_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_1263_n100# a_1215_122# a_1167_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X31 a_1551_n100# a_1503_n188# a_1455_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X32 a_n945_n100# a_n993_n188# a_n1041_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X33 a_n753_n100# a_n801_n188# a_n849_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X34 a_n657_n100# a_n705_122# a_n753_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X35 a_n465_n100# a_n513_122# a_n561_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X36 a_n369_n100# a_n417_n188# a_n465_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X37 a_1167_n100# a_1119_n188# a_1071_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X38 a_1359_n100# a_1311_n188# a_1263_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X39 a_1455_n100# a_1407_122# a_1359_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X40 a_1647_n100# a_1599_122# a_1551_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X41 a_1743_n100# a_1695_n188# a_1647_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X42 a_1935_n100# a_1887_n188# a_1839_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X43 a_n849_n100# a_n897_122# a_n945_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X44 a_1839_n100# a_1791_122# a_1743_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X45 a_15_n100# a_n33_n188# a_n81_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X46 a_n81_n100# a_n129_122# a_n177_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X47 a_111_n100# a_63_122# a_15_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X48 a_n273_n100# a_n321_122# a_n369_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X49 a_n177_n100# a_n225_n188# a_n273_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X50 a_n2865_n100# a_n2913_n188# a_n2957_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X51 a_n2769_n100# a_n2817_122# a_n2865_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X52 a_2127_n100# a_2079_n188# a_2031_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X53 a_2223_n100# a_2175_122# a_2127_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X54 a_2415_n100# a_2367_122# a_2319_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X55 a_2511_n100# a_2463_n188# a_2415_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X56 a_2703_n100# a_2655_n188# a_2607_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X57 a_2319_n100# a_2271_n188# a_2223_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X58 a_2607_n100# a_2559_122# a_2511_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X59 a_2799_n100# a_2751_122# a_2703_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X60 a_2895_n100# a_2847_n188# a_2799_n100# a_n3059_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_4C7XCD a_n573_n491# a_n573_59# a_n703_n621#
X0 a_n573_n491# a_n573_59# a_n703_n621# sky130_fd_pr__res_xhigh_po_5p73 l=590000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_G3ZQK6 a_543_n100# a_7455_n100# a_n609_n100# a_159_n100#
+ a_1695_n100# a_4575_n100# a_3951_122# a_n2001_122# a_2655_n100# a_5535_n100# a_879_122#
+ a_n5793_n100# a_8175_122# a_n7281_n188# a_3615_n100# a_n3873_n100# a_n6753_n100#
+ a_6063_122# a_n2481_n188# a_n5361_n188# a_n8241_n188# a_n6369_n100# a_n7713_n100#
+ a_n273_122# a_n1953_n100# a_n3489_n100# a_n4833_n100# a_n2097_n188# a_n3441_n188#
+ a_n6321_n188# a_n1569_n100# a_n2913_n100# a_n4449_n100# a_n7329_n100# a_n1521_n188#
+ a_n3057_n188# a_n4401_n188# a_n2529_n100# a_n5409_n100# a_1839_122# a_n1137_n188#
+ a_n4017_n188# a_n7569_122# a_n5457_122# a_6591_n100# a_n3345_122# a_n705_n100# a_1791_n100#
+ a_4671_n100# a_7551_n100# a_n1233_122# a_255_n100# a_7167_n100# a_4911_122# a_2751_n100#
+ a_4287_n100# a_5631_n100# a_975_n188# a_2367_n100# a_5247_n100# a_8127_n100# a_7887_n188#
+ a_3711_n100# a_7023_122# a_5967_n188# a_5295_122# a_3327_n100# a_6207_n100# a_n3585_n100#
+ a_n6465_n100# a_6927_n188# a_3183_122# a_1407_n100# a_n7425_n100# a_n1665_n100#
+ a_n4545_n100# a_1071_122# a_n2625_n100# a_n5505_n100# a_n4689_122# a_n6417_122#
+ a_n2577_122# a_n4305_122# a_n801_n100# a_351_n100# a_n417_n100# a_4383_n100# a_7263_n100#
+ a_n7761_122# a_2463_n100# a_5343_n100# a_8223_n100# a_2079_n100# a_6303_n100# a_6255_122#
+ a_n465_122# a_3423_n100# a_n6561_n100# a_n8097_n100# a_4143_122# a_1503_n100# a_3039_n100#
+ a_n3681_n100# a_n1761_n100# a_n3297_n100# a_n4641_n100# a_n6177_n100# a_n7521_n100#
+ a_2031_122# a_1119_n100# a_n6897_n188# a_n1377_n100# a_n2721_n100# a_n4257_n100#
+ a_n5601_n100# a_n7137_n100# a_n5217_n100# a_n4977_n188# a_n7857_n188# a_n2337_n100#
+ a_n5649_122# a_n3537_122# a_n5937_n188# a_n1425_122# a_n513_n100# a_7599_122# a_n129_n100#
+ a_4095_n100# a_783_n188# a_n6993_122# a_7695_n188# a_7215_122# a_5487_122# a_n4881_122#
+ a_2175_n100# a_5055_n100# a_399_n188# a_6015_n100# a_n8193_n100# a_5775_n188# a_5103_122#
+ a_3375_122# a_2895_n188# a_3135_n100# a_n6273_n100# a_1263_122# a_1215_n100# a_n3393_n100#
+ a_6735_n188# a_3855_n188# a_63_n100# a_n1473_n100# a_n4353_n100# a_n7233_n100# a_4815_n188#
+ a_1935_n188# a_n1089_n100# a_n2433_n100# a_n5313_n100# a_n6609_122# a_n2049_n100#
+ a_n2769_122# a_n3009_n100# a_7071_n100# a_n7953_122# a_n225_n100# a_4191_n100# a_6447_122#
+ a_2271_n100# a_5151_n100# a_8031_n100# a_n657_122# a_n945_n188# a_n5841_122# a_4335_122#
+ a_3231_n100# a_6111_n100# a_927_n100# a_3999_n100# a_6879_n100# a_2223_122# a_1311_n100#
+ a_4959_n100# a_7839_n100# a_7791_122# a_5919_n100# a_n1185_n100# a_n4065_n100# a_n4785_n188#
+ a_n7665_n188# a_n2145_n100# a_n5025_n100# a_n3729_122# a_495_122# a_n2865_n188#
+ a_n5745_n188# a_n3105_n100# a_n1617_122# a_111_122# a_n3825_n188# a_n6705_n188#
+ a_n321_n100# a_n1905_n188# a_7407_122# a_5679_122# a_n6801_122# a_3567_122# a_591_n188#
+ a_n2961_122# a_6975_n100# a_5583_n188# a_1455_122# a_n7185_122# a_639_n100# a_7935_n100#
+ a_n6081_n100# a_8079_n188# a_6543_n188# a_5199_n188# a_3663_n188# a_n5073_122# a_1023_n100#
+ a_n1281_n100# a_n4161_n100# a_n7041_n100# a_7503_n188# a_6159_n188# a_4623_n188#
+ a_3279_n188# a_1743_n188# a_207_n188# a_n5121_n100# a_n8001_n100# a_7119_n188# a_4239_n188#
+ a_n2241_n100# a_n5889_n100# a_2703_n188# a_1359_n188# a_n3201_n100# a_2319_n188#
+ a_n3969_n100# a_n6849_n100# a_n7809_n100# a_n4929_n100# a_6639_122# a_n849_122#
+ a_4527_122# a_2799_122# a_n753_n188# a_n3921_122# a_2415_122# a_n369_n188# a_n8145_122#
+ a_6687_n100# a_n33_n100# a_735_n100# a_7983_122# a_n6033_122# a_1887_n100# a_4767_n100#
+ a_7647_n100# a_n2193_122# a_5871_122# a_2847_n100# a_5727_n100# a_3807_n100# a_n5985_n100#
+ a_687_122# a_n4593_n188# a_n7473_n188# a_n6945_n100# a_n1809_122# a_n7089_n188#
+ a_n8387_n274# a_303_122# a_n2673_n188# a_n5553_n188# a_n7905_n100# a_n2289_n188#
+ a_n3633_n188# a_n5169_n188# a_n6513_n188# a_n8049_n188# a_n1713_n188# a_n3249_n188#
+ a_n6129_n188# a_n897_n100# a_3759_122# a_n1329_n188# a_n4209_n188# a_1647_122# a_n7377_122#
+ a_6783_n100# a_5391_n188# a_n5265_122# a_831_n100# a_4863_n100# a_6399_n100# a_7743_n100#
+ a_447_n100# a_1983_n100# a_6831_122# a_6351_n188# a_3471_n188# a_n3153_122# a_1599_n100#
+ a_2943_n100# a_4479_n100# a_5823_n100# a_7359_n100# a_n8285_n100# a_7311_n188# a_3087_n188#
+ a_4431_n188# a_2991_122# a_1551_n188# a_n1041_122# a_2559_n100# a_3903_n100# a_5439_n100#
+ a_4047_n188# a_2511_n188# a_1167_n188# a_3519_n100# a_n5697_n100# a_n3777_n100#
+ a_n6657_n100# a_5007_n188# a_2127_n188# a_n1857_n100# a_n4737_n100# a_n7617_n100#
+ a_n81_122# a_n993_n100# a_n2817_n100# a_4719_122# a_15_n188# a_2607_122# a_n561_n188#
+ a_n4497_122# a_n177_n188# a_n6225_122# a_6495_n100# a_n2385_122# a_n4113_122#
X0 a_3903_n100# a_3855_n188# a_3807_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X1 a_3807_n100# a_3759_122# a_3711_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X2 a_3519_n100# a_3471_n188# a_3423_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X3 a_n6561_n100# a_n6609_122# a_n6657_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X4 a_3999_n100# a_3951_122# a_3903_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X5 a_n6753_n100# a_n6801_122# a_n6849_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X6 a_n6465_n100# a_n6513_n188# a_n6561_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X7 a_6111_n100# a_6063_122# a_6015_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X8 a_n6945_n100# a_n6993_122# a_n7041_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X9 a_n6657_n100# a_n6705_n188# a_n6753_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X10 a_n6369_n100# a_n6417_122# a_n6465_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X11 a_6591_n100# a_6543_n188# a_6495_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X12 a_6303_n100# a_6255_122# a_6207_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X13 a_n6849_n100# a_n6897_n188# a_n6945_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X14 a_6783_n100# a_6735_n188# a_6687_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X15 a_6495_n100# a_6447_122# a_6399_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X16 a_6207_n100# a_6159_n188# a_6111_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X17 a_6975_n100# a_6927_n188# a_6879_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X18 a_6687_n100# a_6639_122# a_6591_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X19 a_6399_n100# a_6351_n188# a_6303_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X20 a_6879_n100# a_6831_122# a_6783_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X21 a_63_n100# a_15_n188# a_n33_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X22 a_n3201_n100# a_n3249_n188# a_n3297_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X23 a_n3681_n100# a_n3729_122# a_n3777_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X24 a_n3393_n100# a_n3441_n188# a_n3489_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X25 a_n3105_n100# a_n3153_122# a_n3201_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X26 a_n3297_n100# a_n3345_122# a_n3393_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X27 a_n3009_n100# a_n3057_n188# a_n3105_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X28 a_n3873_n100# a_n3921_122# a_n3969_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X29 a_n3585_n100# a_n3633_n188# a_n3681_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X30 a_n3777_n100# a_n3825_n188# a_n3873_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X31 a_n3489_n100# a_n3537_122# a_n3585_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X32 a_3231_n100# a_3183_122# a_3135_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X33 a_3135_n100# a_3087_n188# a_3039_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X34 a_3039_n100# a_2991_122# a_2943_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X35 a_n6081_n100# a_n6129_n188# a_n6177_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X36 a_n6273_n100# a_n6321_n188# a_n6369_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X37 a_n5985_n100# a_n6033_122# a_n6081_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X38 a_n6177_n100# a_n6225_122# a_n6273_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X39 a_5823_n100# a_5775_n188# a_5727_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X40 a_6015_n100# a_5967_n188# a_5919_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X41 a_5727_n100# a_5679_122# a_5631_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X42 a_5919_n100# a_5871_122# a_5823_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X43 a_8223_n100# a_8175_122# a_8127_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.1e+11p pd=2.62e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X44 a_8127_n100# a_8079_n188# a_8031_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X45 a_n2241_n100# a_n2289_n188# a_n2337_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X46 a_n2721_n100# a_n2769_122# a_n2817_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X47 a_n2433_n100# a_n2481_n188# a_n2529_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X48 a_n2145_n100# a_n2193_122# a_n2241_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X49 a_n2049_n100# a_n2097_n188# a_n2145_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X50 a_n2913_n100# a_n2961_122# a_n3009_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X51 a_n2625_n100# a_n2673_n188# a_n2721_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X52 a_n2337_n100# a_n2385_122# a_n2433_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X53 a_n2529_n100# a_n2577_122# a_n2625_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X54 a_2271_n100# a_2223_122# a_2175_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X55 a_n2817_n100# a_n2865_n188# a_n2913_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X56 a_2751_n100# a_2703_n188# a_2655_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X57 a_2463_n100# a_2415_122# a_2367_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X58 a_2175_n100# a_2127_n188# a_2079_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X59 a_2079_n100# a_2031_122# a_1983_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X60 a_2943_n100# a_2895_n188# a_2847_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X61 a_2655_n100# a_2607_122# a_2559_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X62 a_2367_n100# a_2319_n188# a_2271_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X63 a_2559_n100# a_2511_n188# a_2463_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X64 a_n5121_n100# a_n5169_n188# a_n5217_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X65 a_2847_n100# a_2799_122# a_2751_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X66 a_n5313_n100# a_n5361_n188# a_n5409_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X67 a_n5025_n100# a_n5073_122# a_n5121_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X68 a_n5601_n100# a_n5649_122# a_n5697_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X69 a_n5793_n100# a_n5841_122# a_n5889_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X70 a_n5505_n100# a_n5553_n188# a_n5601_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X71 a_n5217_n100# a_n5265_122# a_n5313_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X72 a_n5697_n100# a_n5745_n188# a_n5793_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X73 a_n5409_n100# a_n5457_122# a_n5505_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X74 a_5151_n100# a_5103_122# a_5055_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X75 a_5343_n100# a_5295_122# a_5247_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X76 a_5055_n100# a_5007_n188# a_4959_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X77 a_n5889_n100# a_n5937_n188# a_n5985_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X78 a_5631_n100# a_5583_n188# a_5535_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X79 a_5535_n100# a_5487_122# a_5439_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X80 a_5247_n100# a_5199_n188# a_5151_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X81 a_n8001_n100# a_n8049_n188# a_n8097_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X82 a_5439_n100# a_5391_n188# a_5343_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X83 a_1023_n100# a_975_n188# a_927_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X84 a_n8193_n100# a_n8241_n188# a_n8285_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.1e+11p ps=2.62e+06u w=1e+06u l=150000u
X85 a_927_n100# a_879_122# a_831_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X86 a_n8097_n100# a_n8145_122# a_n8193_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X87 a_8031_n100# a_7983_122# a_7935_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X88 a_n1761_n100# a_n1809_122# a_n1857_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X89 a_n1953_n100# a_n2001_122# a_n2049_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X90 a_n1665_n100# a_n1713_n188# a_n1761_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X91 a_n1569_n100# a_n1617_122# a_n1665_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X92 a_1311_n100# a_1263_122# a_1215_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X93 a_n1857_n100# a_n1905_n188# a_n1953_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X94 a_1791_n100# a_1743_n188# a_1695_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X95 a_1503_n100# a_1455_122# a_1407_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X96 a_1215_n100# a_1167_n188# a_1119_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X97 a_1119_n100# a_1071_122# a_1023_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X98 a_1983_n100# a_1935_n188# a_1887_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X99 a_1695_n100# a_1647_122# a_1599_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X100 a_1407_n100# a_1359_n188# a_1311_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X101 a_n4161_n100# a_n4209_n188# a_n4257_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X102 a_1887_n100# a_1839_122# a_1791_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X103 a_1599_n100# a_1551_n188# a_1503_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X104 a_n4065_n100# a_n4113_122# a_n4161_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X105 a_n4641_n100# a_n4689_122# a_n4737_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X106 a_n4353_n100# a_n4401_n188# a_n4449_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X107 a_n4545_n100# a_n4593_n188# a_n4641_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X108 a_n4257_n100# a_n4305_122# a_n4353_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X109 a_n4833_n100# a_n4881_122# a_n4929_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X110 a_n4737_n100# a_n4785_n188# a_n4833_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X111 a_n4449_n100# a_n4497_122# a_n4545_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X112 a_4191_n100# a_4143_122# a_4095_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X113 a_4095_n100# a_4047_n188# a_3999_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X114 a_n33_n100# a_n81_122# a_n129_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X115 a_n4929_n100# a_n4977_n188# a_n5025_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X116 a_4671_n100# a_4623_n188# a_4575_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X117 a_4383_n100# a_4335_122# a_4287_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X118 a_4575_n100# a_4527_122# a_4479_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X119 a_4287_n100# a_4239_n188# a_4191_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X120 a_4863_n100# a_4815_n188# a_4767_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X121 a_n7041_n100# a_n7089_n188# a_n7137_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X122 a_4767_n100# a_4719_122# a_4671_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X123 a_4479_n100# a_4431_n188# a_4383_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X124 a_n7521_n100# a_n7569_122# a_n7617_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X125 a_n7233_n100# a_n7281_n188# a_n7329_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X126 a_4959_n100# a_4911_122# a_4863_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X127 a_351_n100# a_303_122# a_255_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X128 a_n7713_n100# a_n7761_122# a_n7809_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X129 a_n7425_n100# a_n7473_n188# a_n7521_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X130 a_n7137_n100# a_n7185_122# a_n7233_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X131 a_831_n100# a_783_n188# a_735_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X132 a_543_n100# a_495_122# a_447_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X133 a_255_n100# a_207_n188# a_159_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X134 a_n7329_n100# a_n7377_122# a_n7425_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X135 a_7071_n100# a_7023_122# a_6975_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X136 a_n7905_n100# a_n7953_122# a_n8001_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X137 a_n7617_n100# a_n7665_n188# a_n7713_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X138 a_735_n100# a_687_122# a_639_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X139 a_447_n100# a_399_n188# a_351_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X140 a_159_n100# a_111_122# a_63_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X141 a_n7809_n100# a_n7857_n188# a_n7905_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X142 a_7551_n100# a_7503_n188# a_7455_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X143 a_7263_n100# a_7215_122# a_7167_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X144 a_639_n100# a_591_n188# a_543_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X145 a_7743_n100# a_7695_n188# a_7647_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X146 a_7455_n100# a_7407_122# a_7359_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X147 a_7167_n100# a_7119_n188# a_7071_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X148 a_7359_n100# a_7311_n188# a_7263_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X149 a_7935_n100# a_7887_n188# a_7839_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X150 a_7647_n100# a_7599_122# a_7551_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X151 a_n1281_n100# a_n1329_n188# a_n1377_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X152 a_n993_n100# a_n1041_122# a_n1089_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X153 a_7839_n100# a_7791_122# a_7743_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X154 a_n1473_n100# a_n1521_n188# a_n1569_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X155 a_n1185_n100# a_n1233_122# a_n1281_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X156 a_n1377_n100# a_n1425_122# a_n1473_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X157 a_n1089_n100# a_n1137_n188# a_n1185_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X158 a_n321_n100# a_n369_n188# a_n417_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X159 a_n225_n100# a_n273_122# a_n321_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X160 a_n513_n100# a_n561_n188# a_n609_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X161 a_n801_n100# a_n849_122# a_n897_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X162 a_n129_n100# a_n177_n188# a_n225_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X163 a_n417_n100# a_n465_122# a_n513_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X164 a_n705_n100# a_n753_n188# a_n801_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=3.3e+11p pd=2.66e+06u as=0p ps=0u w=1e+06u l=150000u
X165 a_n609_n100# a_n657_122# a_n705_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X166 a_n897_n100# a_n945_n188# a_n993_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X167 a_n3969_n100# a_n4017_n188# a_n4065_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X168 a_3711_n100# a_3663_n188# a_3615_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X169 a_3423_n100# a_3375_122# a_3327_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=3.3e+11p ps=2.66e+06u w=1e+06u l=150000u
X170 a_3615_n100# a_3567_122# a_3519_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
X171 a_3327_n100# a_3279_n188# a_3231_n100# a_n8387_n274# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_HFYJAZ a_15_109# a_n33_n325# a_n33_21# a_n73_n237#
+ a_n73_109# a_15_n237# a_n175_n411#
X0 a_15_n237# a_n33_n325# a_n73_n237# a_n175_n411# sky130_fd_pr__nfet_01v8_lvt ad=1.856e+11p pd=1.86e+06u as=1.856e+11p ps=1.86e+06u w=640000u l=150000u
X1 a_15_109# a_n33_21# a_n73_109# a_n175_n411# sky130_fd_pr__nfet_01v8_lvt ad=1.856e+11p pd=1.86e+06u as=1.856e+11p ps=1.86e+06u w=640000u l=150000u
.ends

.subckt sky130_fd_pr__res_high_po_0p35_C28PVF a_n165_n962# a_n35_n832# a_n35_400#
X0 a_n35_n832# a_n35_400# a_n165_n962# sky130_fd_pr__res_high_po_0p35 l=4e+06u
.ends

.subckt fb vout5p Iref vout5n vin0p vin0n vdd vss
XXM23 vout5n vout5n m1_58226_n6740# vout5n m1_58226_n6740# a_53403_n7310# vout5n vout5n
+ vout5n vout5n m1_58226_n6740# m1_58226_n6740# vout5n m1_58226_n6740# m1_58226_n6740#
+ vout5n vout5n m1_58226_n6740# a_53403_n7310# vout5n vout5n vout5n a_53403_n7310#
+ vss m1_58226_n6740# m1_58226_n6740# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vout5n vout5n m1_58226_n6740# m1_58226_n6740# vout5n m1_58226_n6740# m1_58226_n6740#
+ a_53403_n7310# vout5n vout5n m1_58226_n6740# vout5n vout5n m1_58226_n6740# m1_58226_n6740#
+ vout5n m1_58226_n6740# vout5n a_53403_n7310# vout5n m1_58226_n6740# a_53403_n7310#
+ m1_58226_n6740# vout5n m1_58226_n6740# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# m1_58226_n6740# vout5n m1_58226_n6740# vout5n a_53403_n7310# m1_58226_n6740#
+ m1_58226_n6740# vout5n a_53403_n7310# vout5n vout5n m1_58226_n6740# vout5n vout5n
+ vout5n vout5n vout5n a_53403_n7310# vout5n a_53403_n7310# vout5n vout5n vout5n vout5n
+ vout5n vout5n a_53403_n7310# vout5n a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vout5n a_53403_n7310# vout5n a_53403_n7310# m1_58226_n6740# vout5n a_53403_n7310#
+ m1_58226_n6740# vout5n vout5n vout5n m1_58226_n6740# vout5n vout5n vout5n vout5n
+ m1_58226_n6740# vout5n a_53403_n7310# vout5n a_53403_n7310# vout5n a_53403_n7310#
+ vout5n vout5n vout5n vout5n a_53403_n7310# vout5n m1_58226_n6740# a_53403_n7310#
+ vout5n a_53403_n7310# a_53403_n7310# m1_58226_n6740# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
Xsky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0 m1_58226_n6740# vdd vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXM25 vss vss vss vss vss vss Iref Iref vss vss Iref vss Iref Iref vss vss vss Iref
+ Iref Iref Iref vss vss Iref vss vss vss Iref Iref Iref vss vss vss vss Iref Iref
+ Iref vss vss Iref Iref Iref Iref Iref a_53403_n7310# Iref a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# Iref a_53403_n7310# a_53403_n7310# Iref a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ Iref a_53403_n7310# Iref Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ Iref a_53403_n7310# a_53403_n7310# Iref Iref Iref Iref vss vss vss vss vss Iref
+ vss vss vss vss vss Iref Iref vss vss vss Iref vss vss vss vss vss vss vss vss Iref
+ vss Iref vss vss vss vss vss vss Iref Iref vss Iref Iref Iref Iref a_53403_n7310#
+ Iref a_53403_n7310# a_53403_n7310# Iref Iref Iref Iref Iref Iref a_53403_n7310#
+ a_53403_n7310# Iref a_53403_n7310# a_53403_n7310# Iref Iref Iref Iref a_53403_n7310#
+ a_53403_n7310# Iref a_53403_n7310# a_53403_n7310# Iref Iref a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ Iref a_53403_n7310# Iref a_53403_n7310# vss Iref vss vss Iref vss vss vss Iref Iref
+ Iref Iref vss vss vss vss vss Iref vss vss vss Iref vss vss vss Iref Iref vss vss
+ Iref Iref Iref Iref vss Iref Iref Iref Iref a_53403_n7310# Iref Iref Iref Iref Iref
+ Iref Iref a_53403_n7310# Iref Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ Iref Iref Iref Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ Iref Iref Iref Iref Iref Iref a_53403_n7310# a_53403_n7310# Iref Iref a_53403_n7310#
+ a_53403_n7310# Iref Iref a_53403_n7310# Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# Iref Iref Iref Iref Iref Iref Iref Iref Iref vss vss vss Iref Iref
+ vss vss vss Iref Iref vss vss vss vss Iref Iref Iref vss Iref Iref vss Iref Iref
+ Iref vss Iref Iref Iref Iref Iref Iref Iref Iref a_53403_n7310# Iref Iref Iref Iref
+ Iref a_53403_n7310# Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# Iref Iref Iref Iref a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# a_53403_n7310# vss Iref Iref Iref Iref Iref Iref a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# Iref Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# Iref Iref a_53403_n7310# a_53403_n7310# a_53403_n7310# Iref vss a_53403_n7310#
+ Iref Iref Iref Iref Iref Iref Iref vss Iref Iref sky130_fd_pr__nfet_01v8_lvt_G3ZQK6
Xsky130_fd_pr__nfet_01v8_lvt_HFYJAZ_0 Iref Iref Iref vss vss Iref vss sky130_fd_pr__nfet_01v8_lvt_HFYJAZ
XXR19 vdd m1_48190_n7640# vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
Xsky130_fd_pr__res_high_po_0p35_C28PVF_0 vss m1_48190_n7640# vin0p sky130_fd_pr__res_high_po_0p35_C28PVF
Xsky130_fd_pr__res_high_po_0p35_C28PVF_1 vss m1_58226_n6740# vin0n sky130_fd_pr__res_high_po_0p35_C28PVF
XXM20 vout5p vout5p m1_48190_n7640# vout5p m1_48190_n7640# a_53403_n7310# vout5p vout5p
+ vout5p vout5p m1_48190_n7640# m1_48190_n7640# vout5p m1_48190_n7640# m1_48190_n7640#
+ vout5p vout5p m1_48190_n7640# a_53403_n7310# vout5p vout5p vout5p a_53403_n7310#
+ vss m1_48190_n7640# m1_48190_n7640# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vout5p vout5p m1_48190_n7640# m1_48190_n7640# vout5p m1_48190_n7640# m1_48190_n7640#
+ a_53403_n7310# vout5p vout5p m1_48190_n7640# vout5p vout5p m1_48190_n7640# m1_48190_n7640#
+ vout5p m1_48190_n7640# vout5p a_53403_n7310# vout5p m1_48190_n7640# a_53403_n7310#
+ m1_48190_n7640# vout5p m1_48190_n7640# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# m1_48190_n7640# vout5p m1_48190_n7640# vout5p a_53403_n7310# m1_48190_n7640#
+ m1_48190_n7640# vout5p a_53403_n7310# vout5p vout5p m1_48190_n7640# vout5p vout5p
+ vout5p vout5p vout5p a_53403_n7310# vout5p a_53403_n7310# vout5p vout5p vout5p vout5p
+ vout5p vout5p a_53403_n7310# vout5p a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vout5p a_53403_n7310# vout5p a_53403_n7310# m1_48190_n7640# vout5p a_53403_n7310#
+ m1_48190_n7640# vout5p vout5p vout5p m1_48190_n7640# vout5p vout5p vout5p vout5p
+ m1_48190_n7640# vout5p a_53403_n7310# vout5p a_53403_n7310# vout5p a_53403_n7310#
+ vout5p vout5p vout5p vout5p a_53403_n7310# vout5p m1_48190_n7640# a_53403_n7310#
+ vout5p a_53403_n7310# a_53403_n7310# m1_48190_n7640# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_BSMWRE a_n200_n397# a_200_109# a_n360_n483# a_n200_21#
+ a_200_n309# a_n258_109# a_n258_n309#
X0 a_200_n309# a_n200_n397# a_n258_n309# a_n360_n483# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1 a_200_109# a_n200_21# a_n258_109# a_n360_n483# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_F8HAAN a_n258_1363# a_200_n727# a_n200_n397# a_200_n1145#
+ a_200_109# a_n200_1693# a_n258_n1563# a_n200_857# a_n258_n727# a_n258_527# a_n200_21#
+ a_200_n309# a_n360_n2155# a_200_n1981# a_200_1781# a_n200_n1651# a_200_945# a_n200_1275#
+ a_n200_n2069# a_n258_n1145# a_n200_439# a_n258_109# a_n258_n309# a_n258_1781# a_200_n1563#
+ a_n200_n1233# a_200_1363# a_200_527# a_n258_n1981# a_n200_n815# a_n258_945#
X0 a_200_527# a_n200_439# a_n258_527# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X1 a_200_n309# a_n200_n397# a_n258_n309# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X2 a_200_n1981# a_n200_n2069# a_n258_n1981# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X3 a_200_n1145# a_n200_n1233# a_n258_n1145# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X4 a_200_1363# a_n200_1275# a_n258_1363# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X5 a_200_945# a_n200_857# a_n258_945# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X6 a_200_n727# a_n200_n815# a_n258_n727# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X7 a_200_109# a_n200_21# a_n258_109# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X8 a_200_n1563# a_n200_n1651# a_n258_n1563# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
X9 a_200_1781# a_n200_1693# a_n258_1781# a_n360_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_X3YSY6 w_n246_n319# a_n50_n197# a_50_n100# a_n108_n100#
X0 a_50_n100# a_n50_n197# a_n108_n100# w_n246_n319# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__res_high_po_0p35_ZMQPMJ a_n165_n962# a_n35_n832# a_n35_400#
X0 a_n35_n832# a_n35_400# a_n165_n962# sky130_fd_pr__res_high_po_0p35 l=4e+06u
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_Q3K92U a_n573_n1024# a_n703_n1154# a_n573_592#
X0 a_n573_n1024# a_n573_592# a_n703_n1154# sky130_fd_pr__res_xhigh_po_5p73 l=5.92e+06u
.ends

.subckt sky130_fd_pr__cap_mim_m3_1_L4YDVW c1_n2550_n10450# m3_n2650_n10550#
X0 c1_n2550_n10450# m3_n2650_n10550# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X1 c1_n2550_n10450# m3_n2650_n10550# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X2 c1_n2550_n10450# m3_n2650_n10550# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
X3 c1_n2550_n10450# m3_n2650_n10550# sky130_fd_pr__cap_mim_m3_1 l=2.5e+07u w=2.5e+07u
.ends

.subckt sky130_fd_pr__pfet_01v8_lvt_ER7KZU a_50_1426# a_50_554# a_50_n1190# a_n50_n1723#
+ a_n108_118# a_50_n2062# a_n50_21# a_n108_1426# w_n246_n2281# a_n50_n1287# a_n50_1329#
+ a_n108_n1626# a_n50_n2159# a_50_n754# a_n50_457# a_50_118# a_n108_n754# a_n108_990#
+ a_50_n318# a_n108_n1190# a_n108_n2062# a_n50_n851# a_50_1862# a_50_n1626# a_50_990#
+ a_n108_n318# a_n108_554# a_n108_1862# a_n50_n415# a_n50_1765# a_n50_893#
X0 a_50_1862# a_n50_1765# a_n108_1862# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X1 a_50_n1626# a_n50_n1723# a_n108_n1626# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X2 a_50_n754# a_n50_n851# a_n108_n754# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X3 a_50_n1190# a_n50_n1287# a_n108_n1190# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X4 a_50_118# a_n50_21# a_n108_118# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X5 a_50_n2062# a_n50_n2159# a_n108_n2062# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X6 a_50_554# a_n50_457# a_n108_554# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X7 a_50_990# a_n50_893# a_n108_990# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X8 a_50_1426# a_n50_1329# a_n108_1426# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
X9 a_50_n318# a_n50_n415# a_n108_n318# w_n246_n2281# sky130_fd_pr__pfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=500000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_EA9ZG2 a_25_n100# a_n33_n188# a_n185_n274# a_n83_n100#
X0 a_25_n100# a_n33_n188# a_n83_n100# a_n185_n274# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=250000u
.ends

.subckt cmfb2 vinp vinn vref vc vbcm vdd vss
XXM56 vbcm vss vss vbcm vss m1_n7060_n6640# m1_n7060_n6640# sky130_fd_pr__nfet_01v8_lvt_BSMWRE
XXM57 vc vss vbcm vss vss vbcm vc vbcm vc vc vbcm vss vss vss vss vbcm vss vbcm vbcm
+ vc vbcm vc vc vc vss vbcm vss vss vc vbcm vc sky130_fd_pr__nfet_01v8_lvt_F8HAAN
XXM58 vdd m1_n7220_n6600# m1_n6520_n6580# vdd sky130_fd_pr__pfet_01v8_lvt_X3YSY6
XXM59 vdd m1_n7220_n6600# vdd m1_n7220_n6600# sky130_fd_pr__pfet_01v8_lvt_X3YSY6
XXR34 vss m1_n6520_n6580# m1_n4700_n5960# sky130_fd_pr__res_high_po_0p35_ZMQPMJ
XXR35 vinn vss vcm sky130_fd_pr__res_xhigh_po_5p73_Q3K92U
XXR37 vcm vss vinp sky130_fd_pr__res_xhigh_po_5p73_Q3K92U
XXC4 m1_n4700_n5960# vc sky130_fd_pr__cap_mim_m3_1_L4YDVW
XXM60 vc vc vc m1_n6520_n6580# vdd vc m1_n6520_n6580# vdd vdd m1_n6520_n6580# m1_n6520_n6580#
+ vdd m1_n6520_n6580# vc m1_n6520_n6580# vc vdd vdd vc vdd vdd m1_n6520_n6580# vc
+ vc vc vdd vdd vdd m1_n6520_n6580# m1_n6520_n6580# m1_n6520_n6580# sky130_fd_pr__pfet_01v8_lvt_ER7KZU
XXM54 m1_n7060_n6640# vref vss m1_n7220_n6600# sky130_fd_pr__nfet_01v8_lvt_EA9ZG2
XXM55 m1_n6520_n6580# vcm vss m1_n7060_n6640# sky130_fd_pr__nfet_01v8_lvt_EA9ZG2
.ends

.subckt sky130_fd_pr__res_xhigh_po_5p73_QP6N54 a_n573_150# a_n573_n582# a_n703_n712#
X0 a_n573_n582# a_n573_150# a_n703_n712# sky130_fd_pr__res_xhigh_po_5p73 l=1.5e+06u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_6H2JYD a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt cons_cw voutp vc1 vc2 vinp vinn m1_50970_n6456# m1_47244_n7752# voutn vd22
+ vd21 vss
Xsky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0 vd22 m1_47244_n7752# vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXM23 vinn vinn vd22 vinn vd22 a_53403_n7310# vinn vinn vinn vinn vd22 vd22 vinn vd22
+ vd22 vinn vinn vd22 a_53403_n7310# vinn vinn vinn a_53403_n7310# vss vd22 vd22 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vinn vinn vd22 vd22 vinn vd22 vd22 a_53403_n7310#
+ vinn vinn vd22 vinn vinn vd22 vd22 vinn vd22 vinn a_53403_n7310# vinn vd22 a_53403_n7310#
+ vd22 vinn vd22 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vd22
+ vinn vd22 vinn a_53403_n7310# vd22 vd22 vinn a_53403_n7310# vinn vinn vd22 vinn
+ vinn vinn vinn vinn a_53403_n7310# vinn a_53403_n7310# vinn vinn vinn vinn vinn
+ vinn a_53403_n7310# vinn a_53403_n7310# a_53403_n7310# a_53403_n7310# vinn a_53403_n7310#
+ vinn a_53403_n7310# vd22 vinn a_53403_n7310# vd22 vinn vinn vinn vd22 vinn vinn
+ vinn vinn vd22 vinn a_53403_n7310# vinn a_53403_n7310# vinn a_53403_n7310# vinn
+ vinn vinn vinn a_53403_n7310# vinn vd22 a_53403_n7310# vinn a_53403_n7310# a_53403_n7310#
+ vd22 sky130_fd_pr__nfet_01v8_lvt_FKGFGD
Xsky130_fd_pr__res_xhigh_po_5p73_QP6N54_0 voutn vd22 vss sky130_fd_pr__res_xhigh_po_5p73_QP6N54
XXM24 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# vc2
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vss vc2 vss vss vss vss vc2 vss vss vc2 vss
+ vss vss vc2 vss vss vss vc2 vss vc2 vc2 vc2 vss vss vss vss vc2 vc2 vss vss vss
+ vss vc2 vss vss vc2 vc2 vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 vc2 m1_49981_n5637# vc2 vc2 vc2 vc2 vss vc2 vss vss vc2 vc2 vc2 vc2 vc2 vc2
+ vss vss vc2 vss vss vc2 vc2 vc2 vc2 vss vss vc2 vss vss vc2 vc2 vss vss vss vss
+ vc2 vc2 vss vss vss vc2 vss vc2 vss m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637#
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 vc2 m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637# vc2 vc2
+ vc2 vc2 vss vc2 vc2 vc2 vc2 vc2 vc2 vc2 vss vc2 vc2 vc2 vss vss vss vc2 vc2 vc2
+ vc2 vc2 vss vss vss vss vc2 vc2 vc2 vc2 vc2 vc2 vss vss vc2 vc2 vss vss vc2 vc2
+ vss vc2 vss vss vss vss vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 m1_49981_n5637#
+ vc2 vc2 vss vc2 vc2 vc2 m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 vss vc2
+ vc2 vc2 vc2 vc2 vss vc2 vc2 vss vss vss vss vss vss vc2 vc2 vc2 vc2 vss vss vss
+ vss vss m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vc2 vss vss vss vc2 vc2 vc2 vss vss
+ vss vss vc2 vc2 vss vss vss vc2 m1_49981_n5637# vss vc2 vc2 vc2 vc2 vc2 vc2 vc2
+ m1_49981_n5637# vc2 vc2 sky130_fd_pr__nfet_01v8_lvt_G3ZQK6
XXM25 vss vss vss vss vss vss vc1 vc1 vss vss vc1 vss vc1 vc1 vss vss vss vc1 vc1
+ vc1 vc1 vss vss vc1 vss vss vss vc1 vc1 vc1 vss vss vss vss vc1 vc1 vc1 vss vss
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310#
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vss vss vss vss vss vc1 vss vss vss vss vss vc1 vc1 vss vss vss
+ vc1 vss vss vss vss vss vss vss vss vc1 vss vc1 vss vss vss vss vss vss vc1 vc1
+ vss vc1 vc1 vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1 vc1 vc1
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1
+ vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# vc1 a_53403_n7310# vss vc1 vss
+ vss vc1 vss vss vss vc1 vc1 vc1 vc1 vss vss vss vss vss vc1 vss vss vss vc1 vss
+ vss vss vc1 vc1 vss vss vc1 vc1 vc1 vc1 vss vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310# a_53403_n7310#
+ vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 vc1 vc1 vc1 vc1 vss vss vss vc1 vc1 vss vss vss vc1 vc1 vss
+ vss vss vss vc1 vc1 vc1 vss vc1 vc1 vss vc1 vc1 vc1 vss vc1 vc1 vc1 vc1 vc1 vc1
+ vc1 vc1 a_53403_n7310# vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vss vc1 vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vc1 vss a_53403_n7310# vc1 vc1 vc1 vc1 vc1 vc1 vc1
+ vss vc1 vc1 sky130_fd_pr__nfet_01v8_lvt_G3ZQK6
XXR20 m1_47244_n7752# voutp vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXR21 voutp vd21 vss sky130_fd_pr__res_xhigh_po_5p73_QP6N54
Xsky130_fd_pr__nfet_01v8_lvt_6H2JYD_1 voutn m1_50970_n6456# vd22 vss sky130_fd_pr__nfet_01v8_lvt_6H2JYD
Xsky130_fd_pr__nfet_01v8_lvt_6H2JYD_0 voutp m1_50970_n6456# vd21 vss sky130_fd_pr__nfet_01v8_lvt_6H2JYD
XXR22 voutn m1_47244_n7752# vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXR19 m1_47244_n7752# vd21 vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXM20 vinp vinp vd21 vinp vd21 a_53403_n7310# vinp vinp vinp vinp vd21 vd21 vinp vd21
+ vd21 vinp vinp vd21 a_53403_n7310# vinp vinp vinp a_53403_n7310# vss vd21 vd21 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vinp vinp vd21 vd21 vinp vd21 vd21 a_53403_n7310#
+ vinp vinp vd21 vinp vinp vd21 vd21 vinp vd21 vinp a_53403_n7310# vinp vd21 a_53403_n7310#
+ vd21 vinp vd21 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vd21
+ vinp vd21 vinp a_53403_n7310# vd21 vd21 vinp a_53403_n7310# vinp vinp vd21 vinp
+ vinp vinp vinp vinp a_53403_n7310# vinp a_53403_n7310# vinp vinp vinp vinp vinp
+ vinp a_53403_n7310# vinp a_53403_n7310# a_53403_n7310# a_53403_n7310# vinp a_53403_n7310#
+ vinp a_53403_n7310# vd21 vinp a_53403_n7310# vd21 vinp vinp vinp vd21 vinp vinp
+ vinp vinp vd21 vinp a_53403_n7310# vinp a_53403_n7310# vinp a_53403_n7310# vinp
+ vinp vinp vinp a_53403_n7310# vinp vd21 a_53403_n7310# vinp a_53403_n7310# a_53403_n7310#
+ vd21 sky130_fd_pr__nfet_01v8_lvt_FKGFGD
XXM21 vd21 vd21 m1_49981_n5637# vd21 m1_49981_n5637# voutp vd21 vd21 vd21 vd21 m1_49981_n5637#
+ m1_49981_n5637# vd21 m1_49981_n5637# m1_49981_n5637# vd21 vd21 m1_49981_n5637# voutp
+ vd21 vd21 vd21 voutp vss m1_49981_n5637# m1_49981_n5637# voutp voutp voutp vd21
+ vd21 m1_49981_n5637# m1_49981_n5637# vd21 m1_49981_n5637# m1_49981_n5637# voutp
+ vd21 vd21 m1_49981_n5637# vd21 vd21 m1_49981_n5637# m1_49981_n5637# vd21 m1_49981_n5637#
+ vd21 voutp vd21 m1_49981_n5637# voutp m1_49981_n5637# vd21 m1_49981_n5637# voutp
+ voutp voutp voutp m1_49981_n5637# vd21 m1_49981_n5637# vd21 voutp m1_49981_n5637#
+ m1_49981_n5637# vd21 voutp vd21 vd21 m1_49981_n5637# vd21 vd21 vd21 vd21 vd21 voutp
+ vd21 voutp vd21 vd21 vd21 vd21 vd21 vd21 voutp vd21 voutp voutp voutp vd21 voutp
+ vd21 voutp m1_49981_n5637# vd21 voutp m1_49981_n5637# vd21 vd21 vd21 m1_49981_n5637#
+ vd21 vd21 vd21 vd21 m1_49981_n5637# vd21 voutp vd21 voutp vd21 voutp vd21 vd21 vd21
+ vd21 voutp vd21 m1_49981_n5637# voutp vd21 voutp voutp m1_49981_n5637# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
XXM22 vd22 vd22 m1_49981_n5637# vd22 m1_49981_n5637# voutn vd22 vd22 vd22 vd22 m1_49981_n5637#
+ m1_49981_n5637# vd22 m1_49981_n5637# m1_49981_n5637# vd22 vd22 m1_49981_n5637# voutn
+ vd22 vd22 vd22 voutn vss m1_49981_n5637# m1_49981_n5637# voutn voutn voutn vd22
+ vd22 m1_49981_n5637# m1_49981_n5637# vd22 m1_49981_n5637# m1_49981_n5637# voutn
+ vd22 vd22 m1_49981_n5637# vd22 vd22 m1_49981_n5637# m1_49981_n5637# vd22 m1_49981_n5637#
+ vd22 voutn vd22 m1_49981_n5637# voutn m1_49981_n5637# vd22 m1_49981_n5637# voutn
+ voutn voutn voutn m1_49981_n5637# vd22 m1_49981_n5637# vd22 voutn m1_49981_n5637#
+ m1_49981_n5637# vd22 voutn vd22 vd22 m1_49981_n5637# vd22 vd22 vd22 vd22 vd22 voutn
+ vd22 voutn vd22 vd22 vd22 vd22 vd22 vd22 voutn vd22 voutn voutn voutn vd22 voutn
+ vd22 voutn m1_49981_n5637# vd22 voutn m1_49981_n5637# vd22 vd22 vd22 m1_49981_n5637#
+ vd22 vd22 vd22 vd22 m1_49981_n5637# vd22 voutn vd22 voutn vd22 voutn vd22 vd22 vd22
+ vd22 voutn vd22 m1_49981_n5637# voutn vd22 voutn voutn m1_49981_n5637# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
.ends

.subckt cmfb1 vinn vref vc vbcm vdd vinp vss
XXM56 vbcm vss vss vbcm vss m1_n7060_n6640# m1_n7060_n6640# sky130_fd_pr__nfet_01v8_lvt_BSMWRE
XXM57 vc vss vbcm vss vss vbcm vc vbcm vc vc vbcm vss vss vss vss vbcm vss vbcm vbcm
+ vc vbcm vc vc vc vss vbcm vss vss vc vbcm vc sky130_fd_pr__nfet_01v8_lvt_F8HAAN
XXM58 vdd m1_n7220_n6600# m1_n6520_n6580# vdd sky130_fd_pr__pfet_01v8_lvt_X3YSY6
XXM59 vdd m1_n7220_n6600# vdd m1_n7220_n6600# sky130_fd_pr__pfet_01v8_lvt_X3YSY6
XXR34 vss m1_n6520_n6580# m1_n4700_n5960# sky130_fd_pr__res_high_po_0p35_ZMQPMJ
XXR35 vinn vss vcm sky130_fd_pr__res_xhigh_po_5p73_Q3K92U
XXR37 vcm vss vinp sky130_fd_pr__res_xhigh_po_5p73_Q3K92U
XXC4 m1_n4700_n5960# vc sky130_fd_pr__cap_mim_m3_1_L4YDVW
XXM60 vc vc vc m1_n6520_n6580# vdd vc m1_n6520_n6580# vdd vdd m1_n6520_n6580# m1_n6520_n6580#
+ vdd m1_n6520_n6580# vc m1_n6520_n6580# vc vdd vdd vc vdd vdd m1_n6520_n6580# vc
+ vc vc vdd vdd vdd m1_n6520_n6580# m1_n6520_n6580# m1_n6520_n6580# sky130_fd_pr__pfet_01v8_lvt_ER7KZU
XXM54 m1_n7060_n6640# vref vss m1_n7220_n6600# sky130_fd_pr__nfet_01v8_lvt_EA9ZG2
XXM55 m1_n6520_n6580# vcm vss m1_n7060_n6640# sky130_fd_pr__nfet_01v8_lvt_EA9ZG2
.ends

.subckt stage1 vout1p vout2p vout1n vout2n m1_110_1770# cmfb2_0/vdd vref cmfb2_0/vbcm
+ VSUBS
Xcmfb2_0 vd22 vd21 vref vo21 cmfb2_0/vbcm cmfb2_0/vdd VSUBS cmfb2
Xcons_cw_0 vout2p vo21 vo22 vout1p vout1n m1_110_1770# cmfb2_0/vdd vout2n vd22 vd21
+ VSUBS cons_cw
Xcmfb1_0 vout2p vref vo22 cmfb2_0/vbcm cmfb2_0/vdd vout2n VSUBS cmfb1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_72NHPP a_n33_n1651# a_n73_1363# a_15_1781# a_n33_n815#
+ a_n33_439# a_n33_n2069# a_n33_n397# a_15_109# a_n175_n2155# a_15_n1563# a_n73_n1145#
+ a_n73_n727# a_n73_527# a_15_1363# a_n33_1693# a_n33_n1233# a_n33_21# a_15_945# a_15_n1145#
+ a_n73_n309# a_15_n727# a_n73_109# a_n33_1275# a_n73_n1981# a_n73_1781# a_n33_857#
+ a_15_527# a_15_n1981# a_15_n309# a_n73_n1563# a_n73_945#
X0 a_15_n1145# a_n33_n1233# a_n73_n1145# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1 a_15_1363# a_n33_1275# a_n73_1363# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X2 a_15_n727# a_n33_n815# a_n73_n727# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X3 a_15_527# a_n33_439# a_n73_527# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X4 a_15_n1563# a_n33_n1651# a_n73_n1563# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X5 a_15_1781# a_n33_1693# a_n73_1781# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X6 a_15_945# a_n33_857# a_n73_945# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X7 a_15_n309# a_n33_n397# a_n73_n309# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X8 a_15_109# a_n33_21# a_n73_109# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X9 a_15_n1981# a_n33_n2069# a_n73_n1981# a_n175_n2155# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_8PSHEW a_n33_n216# a_n73_n128# a_15_n128# a_n175_n302#
X0 a_15_n128# a_n33_n216# a_n73_n128# a_n175_n302# sky130_fd_pr__nfet_01v8_lvt ad=3.712e+11p pd=3.14e+06u as=3.712e+11p ps=3.14e+06u w=1.28e+06u l=150000u
.ends

.subckt cons1 voutp vc1 vc2 vinp vinn m1_47244_n7752# voutn vd22 vd21 vss
Xsky130_fd_pr__res_xhigh_po_5p73_4C7XCD_0 vd22 m1_47244_n7752# vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXM23 vinn vinn vd22 vinn vd22 a_53403_n7310# vinn vinn vinn vinn vd22 vd22 vinn vd22
+ vd22 vinn vinn vd22 a_53403_n7310# vinn vinn vinn a_53403_n7310# vss vd22 vd22 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vinn vinn vd22 vd22 vinn vd22 vd22 a_53403_n7310#
+ vinn vinn vd22 vinn vinn vd22 vd22 vinn vd22 vinn a_53403_n7310# vinn vd22 a_53403_n7310#
+ vd22 vinn vd22 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vd22
+ vinn vd22 vinn a_53403_n7310# vd22 vd22 vinn a_53403_n7310# vinn vinn vd22 vinn
+ vinn vinn vinn vinn a_53403_n7310# vinn a_53403_n7310# vinn vinn vinn vinn vinn
+ vinn a_53403_n7310# vinn a_53403_n7310# a_53403_n7310# a_53403_n7310# vinn a_53403_n7310#
+ vinn a_53403_n7310# vd22 vinn a_53403_n7310# vd22 vinn vinn vinn vd22 vinn vinn
+ vinn vinn vd22 vinn a_53403_n7310# vinn a_53403_n7310# vinn a_53403_n7310# vinn
+ vinn vinn vinn a_53403_n7310# vinn vd22 a_53403_n7310# vinn a_53403_n7310# a_53403_n7310#
+ vd22 sky130_fd_pr__nfet_01v8_lvt_FKGFGD
Xsky130_fd_pr__res_xhigh_po_5p73_QP6N54_0 voutn vd22 vss sky130_fd_pr__res_xhigh_po_5p73_QP6N54
XXM24 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# vc2
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vss vc2 vss vss vss vss vc2 vss vss vc2 vss
+ vss vss vc2 vss vss vss vc2 vss vc2 vc2 vc2 vss vss vss vss vc2 vc2 vss vss vss
+ vss vc2 vss vss vc2 vc2 vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 vc2 m1_49981_n5637# vc2 vc2 vc2 vc2 vss vc2 vss vss vc2 vc2 vc2 vc2 vc2 vc2
+ vss vss vc2 vss vss vc2 vc2 vc2 vc2 vss vss vc2 vss vss vc2 vc2 vss vss vss vss
+ vc2 vc2 vss vss vss vc2 vss vc2 vss m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637#
+ vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637#
+ m1_49981_n5637# m1_49981_n5637# vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637#
+ vc2 vc2 m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 vc2 m1_49981_n5637# vc2 vc2
+ vc2 vc2 vss vc2 vc2 vc2 vc2 vc2 vc2 vc2 vss vc2 vc2 vc2 vss vss vss vc2 vc2 vc2
+ vc2 vc2 vss vss vss vss vc2 vc2 vc2 vc2 vc2 vc2 vss vss vc2 vc2 vss vss vc2 vc2
+ vss vc2 vss vss vss vss vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 m1_49981_n5637# m1_49981_n5637#
+ m1_49981_n5637# vc2 vc2 m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2
+ m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# m1_49981_n5637# vc2 vc2 vc2 m1_49981_n5637#
+ vc2 vc2 vss vc2 vc2 vc2 m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vc2 vc2 vc2 vss vc2
+ vc2 vc2 vc2 vc2 vss vc2 vc2 vss vss vss vss vss vss vc2 vc2 vc2 vc2 vss vss vss
+ vss vss m1_49981_n5637# vc2 vc2 vc2 vc2 vc2 vc2 vss vss vss vc2 vc2 vc2 vss vss
+ vss vss vc2 vc2 vss vss vss vc2 m1_49981_n5637# vss vc2 vc2 vc2 vc2 vc2 vc2 vc2
+ m1_49981_n5637# vc2 vc2 sky130_fd_pr__nfet_01v8_lvt_G3ZQK6
XXM25 vss vss vss vss vss vss vc1 vc1 vss vss vc1 vss vc1 vc1 vss vss vss vc1 vc1
+ vc1 vc1 vss vss vc1 vss vss vss vc1 vc1 vc1 vss vss vss vss vc1 vc1 vc1 vss vss
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310#
+ a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310#
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vss vss vss vss vss vc1 vss vss vss vss vss vc1 vc1 vss vss vss
+ vc1 vss vss vss vss vss vss vss vss vc1 vss vc1 vss vss vss vss vss vss vc1 vc1
+ vss vc1 vc1 vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1 vc1 vc1
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1
+ vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# vc1
+ vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vc1 a_53403_n7310# vc1 a_53403_n7310# vss vc1 vss
+ vss vc1 vss vss vss vc1 vc1 vc1 vc1 vss vss vss vss vss vc1 vss vss vss vc1 vss
+ vss vss vc1 vc1 vss vss vc1 vc1 vc1 vc1 vss vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310# a_53403_n7310#
+ vc1 vc1 a_53403_n7310# vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vc1 vc1 vc1 vc1 vc1 vc1 vc1 vc1 vc1 vss vss vss vc1 vc1 vss vss vss vc1 vc1 vss
+ vss vss vss vc1 vc1 vc1 vss vc1 vc1 vss vc1 vc1 vc1 vss vc1 vc1 vc1 vc1 vc1 vc1
+ vc1 vc1 a_53403_n7310# vc1 vc1 vc1 vc1 vc1 a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310#
+ vss vc1 vc1 vc1 vc1 vc1 vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1
+ vc1 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vc1 vc1 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vc1 vss a_53403_n7310# vc1 vc1 vc1 vc1 vc1 vc1 vc1
+ vss vc1 vc1 sky130_fd_pr__nfet_01v8_lvt_G3ZQK6
XXR20 m1_47244_n7752# voutp vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXR21 voutp vd21 vss sky130_fd_pr__res_xhigh_po_5p73_QP6N54
XXR22 voutn m1_47244_n7752# vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXR19 m1_47244_n7752# vd21 vss sky130_fd_pr__res_xhigh_po_5p73_4C7XCD
XXM20 vinp vinp vd21 vinp vd21 a_53403_n7310# vinp vinp vinp vinp vd21 vd21 vinp vd21
+ vd21 vinp vinp vd21 a_53403_n7310# vinp vinp vinp a_53403_n7310# vss vd21 vd21 a_53403_n7310#
+ a_53403_n7310# a_53403_n7310# vinp vinp vd21 vd21 vinp vd21 vd21 a_53403_n7310#
+ vinp vinp vd21 vinp vinp vd21 vd21 vinp vd21 vinp a_53403_n7310# vinp vd21 a_53403_n7310#
+ vd21 vinp vd21 a_53403_n7310# a_53403_n7310# a_53403_n7310# a_53403_n7310# vd21
+ vinp vd21 vinp a_53403_n7310# vd21 vd21 vinp a_53403_n7310# vinp vinp vd21 vinp
+ vinp vinp vinp vinp a_53403_n7310# vinp a_53403_n7310# vinp vinp vinp vinp vinp
+ vinp a_53403_n7310# vinp a_53403_n7310# a_53403_n7310# a_53403_n7310# vinp a_53403_n7310#
+ vinp a_53403_n7310# vd21 vinp a_53403_n7310# vd21 vinp vinp vinp vd21 vinp vinp
+ vinp vinp vd21 vinp a_53403_n7310# vinp a_53403_n7310# vinp a_53403_n7310# vinp
+ vinp vinp vinp a_53403_n7310# vinp vd21 a_53403_n7310# vinp a_53403_n7310# a_53403_n7310#
+ vd21 sky130_fd_pr__nfet_01v8_lvt_FKGFGD
XXM21 vd21 vd21 m1_49981_n5637# vd21 m1_49981_n5637# voutp vd21 vd21 vd21 vd21 m1_49981_n5637#
+ m1_49981_n5637# vd21 m1_49981_n5637# m1_49981_n5637# vd21 vd21 m1_49981_n5637# voutp
+ vd21 vd21 vd21 voutp vss m1_49981_n5637# m1_49981_n5637# voutp voutp voutp vd21
+ vd21 m1_49981_n5637# m1_49981_n5637# vd21 m1_49981_n5637# m1_49981_n5637# voutp
+ vd21 vd21 m1_49981_n5637# vd21 vd21 m1_49981_n5637# m1_49981_n5637# vd21 m1_49981_n5637#
+ vd21 voutp vd21 m1_49981_n5637# voutp m1_49981_n5637# vd21 m1_49981_n5637# voutp
+ voutp voutp voutp m1_49981_n5637# vd21 m1_49981_n5637# vd21 voutp m1_49981_n5637#
+ m1_49981_n5637# vd21 voutp vd21 vd21 m1_49981_n5637# vd21 vd21 vd21 vd21 vd21 voutp
+ vd21 voutp vd21 vd21 vd21 vd21 vd21 vd21 voutp vd21 voutp voutp voutp vd21 voutp
+ vd21 voutp m1_49981_n5637# vd21 voutp m1_49981_n5637# vd21 vd21 vd21 m1_49981_n5637#
+ vd21 vd21 vd21 vd21 m1_49981_n5637# vd21 voutp vd21 voutp vd21 voutp vd21 vd21 vd21
+ vd21 voutp vd21 m1_49981_n5637# voutp vd21 voutp voutp m1_49981_n5637# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
XXM22 vd22 vd22 m1_49981_n5637# vd22 m1_49981_n5637# voutn vd22 vd22 vd22 vd22 m1_49981_n5637#
+ m1_49981_n5637# vd22 m1_49981_n5637# m1_49981_n5637# vd22 vd22 m1_49981_n5637# voutn
+ vd22 vd22 vd22 voutn vss m1_49981_n5637# m1_49981_n5637# voutn voutn voutn vd22
+ vd22 m1_49981_n5637# m1_49981_n5637# vd22 m1_49981_n5637# m1_49981_n5637# voutn
+ vd22 vd22 m1_49981_n5637# vd22 vd22 m1_49981_n5637# m1_49981_n5637# vd22 m1_49981_n5637#
+ vd22 voutn vd22 m1_49981_n5637# voutn m1_49981_n5637# vd22 m1_49981_n5637# voutn
+ voutn voutn voutn m1_49981_n5637# vd22 m1_49981_n5637# vd22 voutn m1_49981_n5637#
+ m1_49981_n5637# vd22 voutn vd22 vd22 m1_49981_n5637# vd22 vd22 vd22 vd22 vd22 voutn
+ vd22 voutn vd22 vd22 vd22 vd22 vd22 vd22 voutn vd22 voutn voutn voutn vd22 voutn
+ vd22 voutn m1_49981_n5637# vd22 voutn m1_49981_n5637# vd22 vd22 vd22 m1_49981_n5637#
+ vd22 vd22 vd22 vd22 m1_49981_n5637# vd22 voutn vd22 voutn vd22 voutn vd22 vd22 vd22
+ vd22 voutn vd22 m1_49981_n5637# voutn vd22 voutn voutn m1_49981_n5637# sky130_fd_pr__nfet_01v8_lvt_FKGFGD
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_L3LEKD a_n258_n100# a_n200_n188# a_n360_n274#
+ a_200_n100#
X0 a_200_n100# a_n200_n188# a_n258_n100# a_n360_n274# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=2e+06u
.ends

.subckt stage0 vout1p vout2p vout1n vout2n vd22 vd21 cmfb2_0/vdd vref cmfb2_0/vbcm
+ VSUBS
Xcmfb2_0 vd22 vd21 vref vo21 cmfb2_0/vbcm cmfb2_0/vdd VSUBS cmfb2
Xcons1_0 vout2p vo21 vo22 vout1p vout1n cmfb2_0/vdd vout2n vd22 vd21 VSUBS cons1
Xsky130_fd_pr__nfet_01v8_lvt_L3LEKD_0 VSUBS cmfb2_0/vbcm VSUBS cmfb2_0/vbcm sky130_fd_pr__nfet_01v8_lvt_L3LEKD
Xcmfb1_0 vout2p vref vo22 cmfb2_0/vbcm cmfb2_0/vdd vout2n VSUBS cmfb1
.ends

.subckt sky130_fd_pr__nfet_01v8_lvt_XA5MKQ a_n33_n1651# a_n73_1363# a_15_1781# a_15_2617#
+ a_n33_2947# a_15_n5325# a_n73_n3235# a_15_n2399# a_n73_3035# a_15_3453# a_n33_3783#
+ a_n33_4619# a_n73_n4071# a_n33_n3323# a_n33_n815# a_n33_439# a_15_2199# a_15_5125#
+ a_n33_5455# a_n33_n2069# a_n33_n397# a_n33_n4995# a_15_109# a_15_n1563# a_n175_n5917#
+ a_n73_n1145# a_n73_n727# a_15_n3235# a_n73_527# a_15_1363# a_n33_1693# a_n33_2529#
+ a_15_n4071# a_n33_n1233# a_n73_n4907# a_15_3035# a_n33_3365# a_n73_3871# a_n73_4707#
+ a_n73_n5743# a_n33_5037# a_n73_5543# a_n33_n5831# a_n73_n4489# a_n33_21# a_n73_4289#
+ a_n33_n4577# a_15_945# a_15_n1145# a_n73_n309# a_15_n727# a_n73_109# a_n33_1275#
+ a_n33_4201# a_15_n4907# a_n73_n2817# a_n73_n1981# a_n73_1781# a_n73_2617# a_n73_n3653#
+ a_n33_n2905# a_15_n5743# a_n73_3453# a_15_3871# a_15_4707# a_n73_n5325# a_15_n4489#
+ a_n33_n3741# a_n73_n2399# a_n33_n5413# a_n33_n2487# a_n33_857# a_n73_2199# a_n73_5125#
+ a_15_5543# a_n33_n4159# a_15_4289# a_15_527# a_n33_2111# a_15_n2817# a_15_n1981#
+ a_15_n309# a_15_n3653# a_n73_n1563# a_n73_945#
X0 a_15_n1145# a_n33_n1233# a_n73_n1145# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X1 a_15_5543# a_n33_5455# a_n73_5543# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X2 a_15_4707# a_n33_4619# a_n73_4707# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X3 a_15_3453# a_n33_3365# a_n73_3453# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X4 a_15_2617# a_n33_2529# a_n73_2617# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X5 a_15_n4489# a_n33_n4577# a_n73_n4489# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X6 a_15_1363# a_n33_1275# a_n73_1363# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X7 a_15_n2399# a_n33_n2487# a_n73_n2399# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X8 a_15_n727# a_n33_n815# a_n73_n727# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X9 a_15_n4907# a_n33_n4995# a_n73_n4907# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X10 a_15_n5743# a_n33_n5831# a_n73_n5743# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X11 a_15_527# a_n33_439# a_n73_527# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X12 a_15_n2817# a_n33_n2905# a_n73_n2817# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X13 a_15_n3653# a_n33_n3741# a_n73_n3653# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X14 a_15_n1563# a_n33_n1651# a_n73_n1563# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X15 a_15_5125# a_n33_5037# a_n73_5125# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X16 a_15_3871# a_n33_3783# a_n73_3871# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X17 a_15_3035# a_n33_2947# a_n73_3035# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X18 a_15_1781# a_n33_1693# a_n73_1781# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X19 a_15_4289# a_n33_4201# a_n73_4289# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X20 a_15_945# a_n33_857# a_n73_945# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X21 a_15_n309# a_n33_n397# a_n73_n309# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X22 a_15_n5325# a_n33_n5413# a_n73_n5325# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X23 a_15_2199# a_n33_2111# a_n73_2199# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X24 a_15_109# a_n33_21# a_n73_109# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X25 a_15_n1981# a_n33_n2069# a_n73_n1981# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X26 a_15_n3235# a_n33_n3323# a_n73_n3235# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
X27 a_15_n4071# a_n33_n4159# a_n73_n4071# a_n175_n5917# sky130_fd_pr__nfet_01v8_lvt ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
.ends

.subckt top vout5p fb_0/vdd fb_0/vout5n vc vin0p vin0n stage0_0/vout1p fb_0/Iref stage0_0/vout1n
+ vref VSUBS
Xfb_0 vout5p fb_0/Iref fb_0/vout5n vin0p vin0n fb_0/vdd VSUBS fb
Xstage1_0 stage1_0/vout1p stage1_1/vout1p stage1_0/vout1n stage1_1/vout1n vc fb_0/vdd
+ vref fb_0/Iref VSUBS stage1
Xstage1_1 stage1_1/vout1p stage1_2/vout1p stage1_1/vout1n stage1_2/vout1n vc fb_0/vdd
+ vref fb_0/Iref VSUBS stage1
Xstage1_2 stage1_2/vout1p stage1_3/vout1p stage1_2/vout1n stage1_3/vout1n vc fb_0/vdd
+ vref fb_0/Iref VSUBS stage1
Xstage1_3 stage1_3/vout1p vout5p stage1_3/vout1n fb_0/vout5n vc fb_0/vdd vref fb_0/Iref
+ VSUBS stage1
Xsky130_fd_pr__nfet_01v8_lvt_72NHPP_0 vin0p m1_5064_n59754# stage0_0/vd21 vin0p vin0p
+ vin0p vin0p stage0_0/vd21 VSUBS stage0_0/vd21 m1_5064_n59754# m1_5064_n59754# m1_5064_n59754#
+ stage0_0/vd21 vin0p vin0p vin0p stage0_0/vd21 stage0_0/vd21 m1_5064_n59754# stage0_0/vd21
+ m1_5064_n59754# vin0p m1_5064_n59754# m1_5064_n59754# vin0p stage0_0/vd21 stage0_0/vd21
+ stage0_0/vd21 m1_5064_n59754# m1_5064_n59754# sky130_fd_pr__nfet_01v8_lvt_72NHPP
Xsky130_fd_pr__nfet_01v8_lvt_8PSHEW_0 fb_0/Iref VSUBS fb_0/Iref VSUBS sky130_fd_pr__nfet_01v8_lvt_8PSHEW
Xsky130_fd_pr__nfet_01v8_lvt_72NHPP_1 vin0n m1_5064_n59754# stage0_0/vd22 vin0n vin0n
+ vin0n vin0n stage0_0/vd22 VSUBS stage0_0/vd22 m1_5064_n59754# m1_5064_n59754# m1_5064_n59754#
+ stage0_0/vd22 vin0n vin0n vin0n stage0_0/vd22 stage0_0/vd22 m1_5064_n59754# stage0_0/vd22
+ m1_5064_n59754# vin0n m1_5064_n59754# m1_5064_n59754# vin0n stage0_0/vd22 stage0_0/vd22
+ stage0_0/vd22 m1_5064_n59754# m1_5064_n59754# sky130_fd_pr__nfet_01v8_lvt_72NHPP
Xstage0_0 stage0_0/vout1p stage1_0/vout1p stage0_0/vout1n stage1_0/vout1n stage0_0/vd22
+ stage0_0/vd21 fb_0/vdd vref fb_0/Iref VSUBS stage0
Xsky130_fd_pr__nfet_01v8_lvt_XA5MKQ_0 fb_0/Iref VSUBS m1_5064_n59754# m1_5064_n59754#
+ fb_0/Iref m1_5064_n59754# VSUBS m1_5064_n59754# VSUBS m1_5064_n59754# fb_0/Iref
+ fb_0/Iref VSUBS fb_0/Iref fb_0/Iref fb_0/Iref m1_5064_n59754# m1_5064_n59754# fb_0/Iref
+ fb_0/Iref fb_0/Iref fb_0/Iref m1_5064_n59754# m1_5064_n59754# VSUBS VSUBS VSUBS
+ m1_5064_n59754# VSUBS m1_5064_n59754# fb_0/Iref fb_0/Iref m1_5064_n59754# fb_0/Iref
+ VSUBS m1_5064_n59754# fb_0/Iref VSUBS VSUBS VSUBS fb_0/Iref VSUBS fb_0/Iref VSUBS
+ fb_0/Iref VSUBS fb_0/Iref m1_5064_n59754# m1_5064_n59754# VSUBS m1_5064_n59754#
+ VSUBS fb_0/Iref fb_0/Iref m1_5064_n59754# VSUBS VSUBS VSUBS VSUBS VSUBS fb_0/Iref
+ m1_5064_n59754# VSUBS m1_5064_n59754# m1_5064_n59754# VSUBS m1_5064_n59754# fb_0/Iref
+ VSUBS fb_0/Iref fb_0/Iref fb_0/Iref VSUBS VSUBS m1_5064_n59754# fb_0/Iref m1_5064_n59754#
+ m1_5064_n59754# fb_0/Iref m1_5064_n59754# m1_5064_n59754# m1_5064_n59754# m1_5064_n59754#
+ VSUBS VSUBS sky130_fd_pr__nfet_01v8_lvt_XA5MKQ
.ends

.subckt VGA_routing top_1/vc top_0/stage0_0/vout1p top_1/fb_0/vout5n top_1/stage0_0/vout1n
+ top_1/vout5p top_0/stage0_0/vout1n top_0/fb_0/Iref top_1/fb_0/Iref top_1/vin0n top_1/stage0_0/vout1p
+ top_1/fb_0/vdd top_1/vin0p top_1/vref VSUBS
Xtop_0 top_1/vout5p top_1/fb_0/vdd top_1/fb_0/vout5n top_1/vc top_1/vin0p top_1/vin0n
+ top_0/stage0_0/vout1p top_0/fb_0/Iref top_0/stage0_0/vout1n top_1/vref VSUBS top
Xtop_1 top_1/vout5p top_1/fb_0/vdd top_1/fb_0/vout5n top_1/vc top_1/vin0p top_1/vin0n
+ top_1/stage0_0/vout1p top_1/fb_0/Iref top_1/stage0_0/vout1n top_1/vref VSUBS top
.ends

.subckt user_analog_project_wrapper gpio_analog[0] gpio_analog[10] gpio_analog[11]
+ gpio_analog[12] gpio_analog[13] gpio_analog[14] gpio_analog[15] gpio_analog[16]
+ gpio_analog[17] gpio_analog[1] gpio_analog[2] gpio_analog[3] gpio_analog[4] gpio_analog[5]
+ gpio_analog[6] gpio_analog[7] gpio_analog[8] gpio_analog[9] gpio_noesd[0] gpio_noesd[10]
+ gpio_noesd[11] gpio_noesd[12] gpio_noesd[13] gpio_noesd[14] gpio_noesd[15] gpio_noesd[16]
+ gpio_noesd[17] gpio_noesd[1] gpio_noesd[2] gpio_noesd[3] gpio_noesd[4] gpio_noesd[5]
+ gpio_noesd[6] gpio_noesd[7] gpio_noesd[8] gpio_noesd[9] io_analog[0] io_analog[1]
+ io_analog[2] io_analog[3] io_analog[6] io_analog[7] io_analog[8] io_analog[9] io_analog[4]
+ io_analog[5] io_clamp_high[0] io_clamp_high[1] io_clamp_high[2] io_clamp_low[0]
+ io_clamp_low[1] io_clamp_low[2] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13]
+ io_in[14] io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21]
+ io_in[22] io_in[23] io_in[24] io_in[25] io_in[26] io_in[2] io_in[3] io_in[4] io_in[5]
+ io_in[6] io_in[7] io_in[8] io_in[9] io_in_3v3[0] io_in_3v3[10] io_in_3v3[11] io_in_3v3[12]
+ io_in_3v3[13] io_in_3v3[14] io_in_3v3[15] io_in_3v3[16] io_in_3v3[17] io_in_3v3[18]
+ io_in_3v3[19] io_in_3v3[1] io_in_3v3[20] io_in_3v3[21] io_in_3v3[22] io_in_3v3[23]
+ io_in_3v3[24] io_in_3v3[25] io_in_3v3[26] io_in_3v3[2] io_in_3v3[3] io_in_3v3[4]
+ io_in_3v3[5] io_in_3v3[6] io_in_3v3[7] io_in_3v3[8] io_in_3v3[9] io_oeb[0] io_oeb[10]
+ io_oeb[11] io_oeb[12] io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18]
+ io_oeb[19] io_oeb[1] io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25]
+ io_oeb[26] io_oeb[2] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7] io_oeb[8]
+ io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14] io_out[15]
+ io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21] io_out[22]
+ io_out[23] io_out[24] io_out[25] io_out[26] io_out[2] io_out[3] io_out[4] io_out[5]
+ io_out[6] io_out[7] io_out[8] io_out[9] la_data_in[0] la_data_in[100] la_data_in[101]
+ la_data_in[102] la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106]
+ la_data_in[107] la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111]
+ la_data_in[112] la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116]
+ la_data_in[117] la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121]
+ la_data_in[122] la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126]
+ la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16]
+ la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21]
+ la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27]
+ la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32]
+ la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38]
+ la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43]
+ la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49]
+ la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54]
+ la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5]
+ la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65]
+ la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70]
+ la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76]
+ la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81]
+ la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87]
+ la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92]
+ la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98]
+ la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] user_clock2 user_irq[0] user_irq[1] user_irq[2]
+ vccd1 vccd2 vdda1 vdda2 vssa1 vssa2 vssd1 vssd2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i io_analog[10]
XVCO_0 REF CTRL5 io_in[18] io_analog[10] io_in[17] vdda2 io_analog[8] io_in[16] io_analog[9]
+ io_in_3v3[15] vssa2 VCO
XVCO_1 REF2 CTRL5 io_in[18] io_analog[10] io_in[17] vdda2 txinb io_in[16] txina io_in_3v3[15]
+ vssa2 VCO
XTX_line_0 txinb txina vssa2 TX_line
XBGR_lvs_0 REF2 REF io_analog[7] gpio_analog[7] io_analog[6] BGR_lvs_0/Iout3 BGR_lvs_0/Iout4
+ BGR_lvs_0/Iout5 BGR_lvs_0/Iout6 vccd2 vssa2 BGR_lvs
XVGA_routing_0 io_in[13] txina io_analog[2] io_analog[5] io_analog[3] txinb BGR_lvs_0/Iout4
+ BGR_lvs_0/Iout3 io_analog[1] io_analog[4] vccd1 io_analog[0] io_analog[6] vssa2
+ VGA_routing
.ends

