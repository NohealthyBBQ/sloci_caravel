magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect 14349 524 14447 776
<< ndiff >>
rect 14375 550 14421 750
<< locali >>
rect 12675 1830 13610 1870
rect 10060 880 10095 1110
rect 12665 1070 13615 1075
rect 11900 925 11935 1070
rect 12055 925 12090 1070
rect 11900 885 12090 925
rect 12665 1035 13630 1070
rect 12665 930 12705 1035
rect 13595 930 13630 1035
rect 12665 890 13630 930
rect 15745 920 15780 1075
rect 15895 920 15930 1070
rect 15745 890 15930 920
rect 17960 890 17995 1140
rect 12665 885 12705 890
rect 15745 885 15925 890
rect 9755 230 9795 420
rect 11905 235 11945 425
rect 12050 230 12090 420
rect 12690 415 13625 420
rect 12665 405 13625 415
rect 12665 380 13635 405
rect 12665 265 12705 380
rect 13600 265 13635 380
rect 12665 225 13635 265
rect 15735 230 15770 410
rect 15910 230 15945 410
rect 21885 225 21920 415
rect 11905 -250 12090 -245
rect 10055 -430 10095 -250
rect 11905 -285 12095 -250
rect 11905 -430 11945 -285
rect 12055 -430 12095 -285
rect 12660 -260 13625 -250
rect 15740 -255 15775 -245
rect 15895 -255 15930 -245
rect 12660 -290 13630 -260
rect 12660 -400 12700 -290
rect 13595 -400 13630 -290
rect 12660 -430 13630 -400
rect 15740 -290 15930 -255
rect 15740 -425 15775 -290
rect 15895 -425 15930 -290
rect 12680 -440 13630 -430
rect 17965 -435 18005 -250
rect 12675 -1220 13610 -1180
<< metal1 >>
rect 13740 2273 14120 2280
rect 10210 1705 10605 1720
rect 10210 1205 10221 1705
rect 10593 1205 10605 1705
rect 10210 1190 10605 1205
rect 12140 1702 12590 1735
rect 12140 1202 12186 1702
rect 12558 1202 12590 1702
rect 12140 1165 12590 1202
rect 13740 1197 13744 2273
rect 14116 1197 14120 2273
rect 13740 1190 14120 1197
rect 17435 2273 17870 2310
rect 17435 1197 17461 2273
rect 17833 1197 17870 2273
rect 17435 1165 17870 1197
rect 13515 848 13590 860
rect 9900 780 11975 830
rect 12190 780 12740 830
rect 13515 796 13526 848
rect 13578 835 13590 848
rect 13578 796 15675 835
rect 13515 785 15675 796
rect 9860 625 9910 750
rect 9945 738 10020 750
rect 9945 686 9956 738
rect 10008 686 10020 738
rect 9945 675 10020 686
rect 9850 613 9925 625
rect 9850 561 9861 613
rect 9913 561 9925 613
rect 9850 550 9925 561
rect 9960 550 10010 675
rect 10050 625 10100 750
rect 10140 738 10215 750
rect 10140 686 10151 738
rect 10203 686 10215 738
rect 10140 675 10215 686
rect 10040 613 10115 625
rect 10040 561 10051 613
rect 10103 561 10115 613
rect 10040 550 10115 561
rect 10150 550 10200 675
rect 10250 625 10300 750
rect 10330 738 10405 750
rect 10330 686 10341 738
rect 10393 686 10405 738
rect 10330 675 10405 686
rect 10230 613 10305 625
rect 10230 561 10241 613
rect 10293 561 10305 613
rect 10230 550 10305 561
rect 10340 550 10390 675
rect 10440 625 10490 750
rect 10520 738 10595 750
rect 10520 686 10531 738
rect 10583 686 10595 738
rect 10520 675 10595 686
rect 10420 613 10495 625
rect 10420 561 10431 613
rect 10483 561 10495 613
rect 10420 550 10495 561
rect 10530 550 10580 675
rect 10630 625 10680 750
rect 10710 738 10785 750
rect 10710 686 10721 738
rect 10773 686 10785 738
rect 10710 675 10785 686
rect 10620 613 10695 625
rect 10620 561 10631 613
rect 10683 561 10695 613
rect 10620 550 10695 561
rect 10730 550 10780 675
rect 10820 625 10870 750
rect 10900 738 10975 750
rect 10900 686 10911 738
rect 10963 686 10975 738
rect 10900 675 10975 686
rect 10810 613 10885 625
rect 10810 561 10821 613
rect 10873 561 10885 613
rect 10810 550 10885 561
rect 10920 550 10970 675
rect 11010 625 11060 750
rect 11095 738 11170 750
rect 11095 686 11106 738
rect 11158 686 11170 738
rect 11095 675 11170 686
rect 11005 613 11080 625
rect 11005 561 11016 613
rect 11068 561 11080 613
rect 11005 550 11080 561
rect 11110 550 11160 675
rect 11210 625 11260 750
rect 11290 738 11365 750
rect 11290 686 11301 738
rect 11353 686 11365 738
rect 11290 675 11365 686
rect 11195 613 11270 625
rect 11195 561 11206 613
rect 11258 561 11270 613
rect 11195 550 11270 561
rect 11300 550 11350 675
rect 11400 625 11450 750
rect 11480 738 11555 750
rect 11480 686 11491 738
rect 11543 686 11555 738
rect 11480 675 11555 686
rect 11385 613 11460 625
rect 11385 561 11396 613
rect 11448 561 11460 613
rect 11385 550 11460 561
rect 11490 550 11540 675
rect 11590 625 11640 750
rect 11675 738 11750 750
rect 11675 686 11686 738
rect 11738 686 11750 738
rect 11675 675 11750 686
rect 11580 613 11655 625
rect 11580 561 11591 613
rect 11643 561 11655 613
rect 11580 550 11655 561
rect 11690 550 11740 675
rect 11780 625 11830 750
rect 11770 613 11845 625
rect 11770 561 11781 613
rect 11833 561 11845 613
rect 11770 550 11845 561
rect 11925 520 11975 780
rect 12165 625 12215 750
rect 12245 738 12320 750
rect 12245 686 12256 738
rect 12308 686 12320 738
rect 12245 675 12320 686
rect 12150 613 12225 625
rect 12150 561 12161 613
rect 12213 561 12225 613
rect 12150 550 12225 561
rect 12255 550 12306 675
rect 12350 625 12401 750
rect 12435 738 12510 750
rect 12435 686 12446 738
rect 12498 686 12510 738
rect 12435 675 12510 686
rect 12340 613 12415 625
rect 12340 561 12351 613
rect 12403 561 12415 613
rect 12340 550 12415 561
rect 12450 550 12501 675
rect 12545 625 12596 750
rect 12535 613 12610 625
rect 12535 561 12546 613
rect 12598 561 12610 613
rect 12535 550 12610 561
rect 12685 520 12740 780
rect 13535 520 13585 785
rect 15855 780 21775 830
rect 13785 738 13860 750
rect 13785 686 13796 738
rect 13848 686 13860 738
rect 13785 675 13860 686
rect 13705 625 13750 670
rect 13690 613 13765 625
rect 13690 561 13701 613
rect 13753 561 13765 613
rect 13690 550 13765 561
rect 13800 550 13846 675
rect 13895 625 13941 750
rect 13975 738 14050 750
rect 13975 686 13986 738
rect 14038 686 14050 738
rect 13975 675 14050 686
rect 13880 613 13955 625
rect 13880 561 13891 613
rect 13943 561 13955 613
rect 13880 550 13955 561
rect 13990 550 14036 675
rect 14085 625 14131 750
rect 14170 738 14245 750
rect 14170 686 14181 738
rect 14233 686 14245 738
rect 14170 675 14245 686
rect 14075 613 14150 625
rect 14075 561 14086 613
rect 14138 561 14150 613
rect 14075 550 14150 561
rect 14185 550 14231 675
rect 14280 625 14326 750
rect 14360 738 14435 750
rect 14360 686 14371 738
rect 14423 686 14435 738
rect 14360 675 14435 686
rect 14265 613 14340 625
rect 14265 561 14276 613
rect 14328 561 14340 613
rect 14265 550 14340 561
rect 14375 550 14421 675
rect 14470 625 14516 750
rect 14550 738 14625 750
rect 14550 686 14561 738
rect 14613 686 14625 738
rect 14550 675 14625 686
rect 14460 613 14535 625
rect 14460 561 14471 613
rect 14523 561 14535 613
rect 14460 550 14535 561
rect 14565 550 14611 675
rect 14665 625 14711 750
rect 14745 738 14820 750
rect 14745 686 14756 738
rect 14808 686 14820 738
rect 14745 675 14820 686
rect 14645 613 14720 625
rect 14645 561 14656 613
rect 14708 561 14720 613
rect 14645 550 14720 561
rect 14760 550 14806 675
rect 14855 625 14901 750
rect 14935 738 15010 750
rect 14935 686 14946 738
rect 14998 686 15010 738
rect 14935 675 15010 686
rect 14840 613 14915 625
rect 14840 561 14851 613
rect 14903 561 14915 613
rect 14840 550 14915 561
rect 14950 550 14996 675
rect 15050 625 15096 750
rect 15130 738 15205 750
rect 15130 686 15141 738
rect 15193 686 15205 738
rect 15130 675 15205 686
rect 15030 613 15105 625
rect 15030 561 15041 613
rect 15093 561 15105 613
rect 15030 550 15105 561
rect 15145 550 15191 675
rect 15240 625 15286 750
rect 15320 738 15395 750
rect 15320 686 15331 738
rect 15383 686 15395 738
rect 15320 675 15395 686
rect 15225 613 15300 625
rect 15225 561 15236 613
rect 15288 561 15300 613
rect 15225 550 15300 561
rect 15335 550 15381 675
rect 15430 625 15476 750
rect 15510 738 15585 750
rect 15510 686 15521 738
rect 15573 686 15585 738
rect 15510 675 15585 686
rect 15415 613 15490 625
rect 15415 561 15426 613
rect 15478 561 15490 613
rect 15415 550 15490 561
rect 15525 550 15571 675
rect 15625 625 15671 750
rect 15610 613 15685 625
rect 15610 561 15621 613
rect 15673 561 15685 613
rect 15610 550 15685 561
rect 9990 470 11975 520
rect 12295 470 13415 520
rect 13535 470 15625 520
rect 15855 515 15905 780
rect 16005 625 16050 750
rect 16085 738 16160 750
rect 16085 686 16096 738
rect 16148 686 16160 738
rect 16085 675 16160 686
rect 15985 613 16060 625
rect 15985 561 15996 613
rect 16048 561 16060 613
rect 15985 550 16060 561
rect 16100 550 16145 675
rect 16195 625 16240 750
rect 16275 738 16350 750
rect 16275 686 16286 738
rect 16338 686 16350 738
rect 16275 675 16350 686
rect 16175 613 16250 625
rect 16175 561 16186 613
rect 16238 561 16250 613
rect 16175 550 16250 561
rect 16290 550 16335 675
rect 16385 625 16430 750
rect 16470 738 16545 750
rect 16470 686 16481 738
rect 16533 686 16545 738
rect 16470 675 16545 686
rect 16370 613 16445 625
rect 16370 561 16381 613
rect 16433 561 16445 613
rect 16370 550 16445 561
rect 16485 550 16530 675
rect 16580 625 16625 750
rect 16660 738 16735 750
rect 16660 686 16671 738
rect 16723 686 16735 738
rect 16660 675 16735 686
rect 16565 613 16640 625
rect 16565 561 16576 613
rect 16628 561 16640 613
rect 16565 550 16640 561
rect 16675 550 16720 675
rect 16770 625 16815 750
rect 16855 738 16930 750
rect 16855 686 16866 738
rect 16918 686 16930 738
rect 16855 675 16930 686
rect 16755 613 16830 625
rect 16755 561 16766 613
rect 16818 561 16830 613
rect 16755 550 16830 561
rect 16870 550 16915 675
rect 16965 625 17010 750
rect 17040 738 17115 750
rect 17040 686 17051 738
rect 17103 686 17115 738
rect 17040 675 17115 686
rect 16950 613 17025 625
rect 16950 561 16961 613
rect 17013 561 17025 613
rect 16950 550 17025 561
rect 17060 550 17105 675
rect 17155 625 17200 750
rect 17240 738 17315 750
rect 17240 686 17251 738
rect 17303 686 17315 738
rect 17240 675 17315 686
rect 17140 613 17215 625
rect 17140 561 17151 613
rect 17203 561 17215 613
rect 17140 550 17215 561
rect 17250 550 17295 675
rect 17350 625 17395 750
rect 17425 738 17500 750
rect 17425 686 17436 738
rect 17488 686 17500 738
rect 17425 675 17500 686
rect 17335 613 17410 625
rect 17335 561 17346 613
rect 17398 561 17410 613
rect 17335 550 17410 561
rect 17445 550 17490 675
rect 17540 625 17585 750
rect 17620 738 17695 750
rect 17620 686 17631 738
rect 17683 686 17695 738
rect 17620 675 17695 686
rect 17525 613 17600 625
rect 17525 561 17536 613
rect 17588 561 17600 613
rect 17525 550 17600 561
rect 17635 550 17680 675
rect 17735 625 17780 750
rect 17815 738 17890 750
rect 17815 686 17826 738
rect 17878 686 17890 738
rect 17815 675 17890 686
rect 17715 613 17790 625
rect 17715 561 17726 613
rect 17778 561 17790 613
rect 17715 550 17790 561
rect 17830 550 17875 675
rect 17925 625 17970 750
rect 18000 738 18075 750
rect 18000 686 18011 738
rect 18063 686 18075 738
rect 18000 675 18075 686
rect 17910 613 17985 625
rect 17910 561 17921 613
rect 17973 561 17985 613
rect 17910 550 17985 561
rect 18020 550 18065 675
rect 18115 625 18160 750
rect 18195 738 18270 750
rect 18195 686 18206 738
rect 18258 686 18270 738
rect 18195 675 18270 686
rect 18100 613 18175 625
rect 18100 561 18111 613
rect 18163 561 18175 613
rect 18100 550 18175 561
rect 18210 550 18255 675
rect 18310 625 18355 750
rect 18385 738 18460 750
rect 18385 686 18396 738
rect 18448 686 18460 738
rect 18385 675 18460 686
rect 18295 613 18370 625
rect 18295 561 18306 613
rect 18358 561 18370 613
rect 18295 550 18370 561
rect 18405 550 18450 675
rect 18500 625 18545 750
rect 18580 738 18655 750
rect 18580 686 18591 738
rect 18643 686 18655 738
rect 18580 675 18655 686
rect 18485 613 18560 625
rect 18485 561 18496 613
rect 18548 561 18560 613
rect 18485 550 18560 561
rect 18595 550 18640 675
rect 18690 625 18735 750
rect 18770 738 18845 750
rect 18770 686 18781 738
rect 18833 686 18845 738
rect 18770 675 18845 686
rect 18675 613 18750 625
rect 18675 561 18686 613
rect 18738 561 18750 613
rect 18675 550 18750 561
rect 18790 550 18835 675
rect 18885 625 18930 750
rect 18965 738 19040 750
rect 18965 686 18976 738
rect 19028 686 19040 738
rect 18965 675 19040 686
rect 18870 613 18945 625
rect 18870 561 18881 613
rect 18933 561 18945 613
rect 18870 550 18945 561
rect 18980 550 19025 675
rect 19075 625 19120 750
rect 19155 738 19230 750
rect 19155 686 19166 738
rect 19218 686 19230 738
rect 19155 675 19230 686
rect 19060 613 19135 625
rect 19060 561 19071 613
rect 19123 561 19135 613
rect 19060 550 19135 561
rect 19170 550 19215 675
rect 19270 625 19315 750
rect 19350 738 19425 750
rect 19350 686 19361 738
rect 19413 686 19425 738
rect 19350 675 19425 686
rect 19255 613 19330 625
rect 19255 561 19266 613
rect 19318 561 19330 613
rect 19255 550 19330 561
rect 19365 550 19410 675
rect 19460 625 19505 750
rect 19540 738 19615 750
rect 19540 686 19551 738
rect 19603 686 19615 738
rect 19540 675 19615 686
rect 19445 613 19520 625
rect 19445 561 19456 613
rect 19508 561 19520 613
rect 19445 550 19520 561
rect 19555 550 19600 675
rect 19650 625 19695 750
rect 19735 738 19810 750
rect 19735 686 19746 738
rect 19798 686 19810 738
rect 19735 675 19810 686
rect 19635 613 19710 625
rect 19635 561 19646 613
rect 19698 561 19710 613
rect 19635 550 19710 561
rect 19750 550 19795 675
rect 19845 625 19890 750
rect 19925 738 20000 750
rect 19925 686 19936 738
rect 19988 686 20000 738
rect 19925 675 20000 686
rect 19830 613 19905 625
rect 19830 561 19841 613
rect 19893 561 19905 613
rect 19830 550 19905 561
rect 19940 550 19985 675
rect 20035 625 20080 750
rect 20115 738 20190 750
rect 20115 686 20126 738
rect 20178 686 20190 738
rect 20115 675 20190 686
rect 20020 613 20095 625
rect 20020 561 20031 613
rect 20083 561 20095 613
rect 20020 550 20095 561
rect 20135 550 20180 675
rect 20230 625 20275 750
rect 20310 738 20385 750
rect 20310 686 20321 738
rect 20373 686 20385 738
rect 20310 675 20385 686
rect 20215 613 20290 625
rect 20215 561 20226 613
rect 20278 561 20290 613
rect 20215 550 20290 561
rect 20325 550 20370 675
rect 20420 625 20465 750
rect 20500 738 20575 750
rect 20500 686 20511 738
rect 20563 686 20575 738
rect 20500 675 20575 686
rect 20405 613 20480 625
rect 20405 561 20416 613
rect 20468 561 20480 613
rect 20405 550 20480 561
rect 20515 550 20560 675
rect 20610 625 20655 750
rect 20695 738 20770 750
rect 20695 686 20706 738
rect 20758 686 20770 738
rect 20695 675 20770 686
rect 20600 613 20675 625
rect 20600 561 20611 613
rect 20663 561 20675 613
rect 20600 550 20675 561
rect 20710 550 20755 675
rect 20805 625 20850 750
rect 20885 738 20960 750
rect 20885 686 20896 738
rect 20948 686 20960 738
rect 20885 675 20960 686
rect 20790 613 20865 625
rect 20790 561 20801 613
rect 20853 561 20865 613
rect 20790 550 20865 561
rect 20900 550 20945 675
rect 20995 625 21040 750
rect 21075 738 21150 750
rect 21075 686 21086 738
rect 21138 686 21150 738
rect 21075 675 21150 686
rect 20980 613 21055 625
rect 20980 561 20991 613
rect 21043 561 21055 613
rect 20980 550 21055 561
rect 21090 550 21135 675
rect 21190 625 21235 750
rect 21270 738 21345 750
rect 21270 686 21281 738
rect 21333 686 21345 738
rect 21270 675 21345 686
rect 21175 613 21250 625
rect 21175 561 21186 613
rect 21238 561 21250 613
rect 21175 550 21250 561
rect 21285 550 21330 675
rect 21380 625 21425 750
rect 21460 738 21535 750
rect 21460 686 21471 738
rect 21523 686 21535 738
rect 21460 675 21535 686
rect 21365 613 21440 625
rect 21365 561 21376 613
rect 21428 561 21440 613
rect 21365 550 21440 561
rect 21475 550 21520 675
rect 21570 625 21615 750
rect 21650 738 21725 750
rect 21650 686 21661 738
rect 21713 686 21725 738
rect 21650 675 21725 686
rect 21555 613 21630 625
rect 21555 561 21566 613
rect 21618 561 21630 613
rect 21555 550 21630 561
rect 21670 550 21715 675
rect 21765 625 21810 750
rect 21750 613 21825 625
rect 21750 561 21761 613
rect 21813 561 21825 613
rect 21750 550 21825 561
rect 11925 170 11975 470
rect 9990 120 11975 170
rect 12290 125 12955 175
rect 12295 120 12955 125
rect 9850 78 9925 90
rect 9850 26 9861 78
rect 9913 26 9925 78
rect 9850 15 9925 26
rect 9860 -110 9910 15
rect 9960 -35 10010 90
rect 10040 78 10115 90
rect 10040 26 10051 78
rect 10103 26 10115 78
rect 10040 15 10115 26
rect 9945 -47 10020 -35
rect 9945 -99 9956 -47
rect 10008 -99 10020 -47
rect 9945 -110 10020 -99
rect 10050 -110 10102 15
rect 10150 -35 10200 90
rect 10230 78 10305 90
rect 10230 26 10241 78
rect 10293 26 10305 78
rect 10230 15 10305 26
rect 10140 -47 10215 -35
rect 10140 -99 10151 -47
rect 10203 -99 10215 -47
rect 10140 -110 10215 -99
rect 10248 -110 10300 15
rect 10340 -35 10390 90
rect 10420 78 10495 90
rect 10420 26 10431 78
rect 10483 26 10495 78
rect 10420 15 10495 26
rect 10330 -47 10405 -35
rect 10330 -99 10341 -47
rect 10393 -99 10405 -47
rect 10330 -110 10405 -99
rect 10440 -110 10490 15
rect 10530 -35 10582 90
rect 10620 78 10695 90
rect 10620 26 10631 78
rect 10683 26 10695 78
rect 10620 15 10695 26
rect 10520 -47 10595 -35
rect 10520 -99 10531 -47
rect 10583 -99 10595 -47
rect 10520 -110 10595 -99
rect 10630 -110 10680 15
rect 10728 -35 10780 90
rect 10810 78 10885 90
rect 10810 26 10821 78
rect 10873 26 10885 78
rect 10810 15 10885 26
rect 10710 -47 10785 -35
rect 10710 -99 10721 -47
rect 10773 -99 10785 -47
rect 10710 -110 10785 -99
rect 10820 -110 10870 15
rect 10920 -35 10970 90
rect 11005 78 11080 90
rect 11005 26 11016 78
rect 11068 26 11080 78
rect 11005 15 11080 26
rect 10900 -47 10975 -35
rect 10900 -99 10911 -47
rect 10963 -99 10975 -47
rect 10900 -110 10975 -99
rect 11010 -110 11062 15
rect 11110 -35 11160 90
rect 11195 78 11270 90
rect 11195 26 11206 78
rect 11258 26 11270 78
rect 11195 15 11270 26
rect 11095 -47 11170 -35
rect 11095 -99 11106 -47
rect 11158 -99 11170 -47
rect 11095 -110 11170 -99
rect 11208 -110 11260 15
rect 11300 -35 11350 90
rect 11385 78 11460 90
rect 11385 26 11396 78
rect 11448 26 11460 78
rect 11385 15 11460 26
rect 11290 -47 11365 -35
rect 11290 -99 11301 -47
rect 11353 -99 11365 -47
rect 11290 -110 11365 -99
rect 11400 -110 11450 15
rect 11490 -35 11542 90
rect 11580 78 11655 90
rect 11580 26 11591 78
rect 11643 26 11655 78
rect 11580 15 11655 26
rect 11480 -47 11555 -35
rect 11480 -99 11491 -47
rect 11543 -99 11555 -47
rect 11480 -110 11555 -99
rect 11590 -110 11640 15
rect 11688 -35 11740 90
rect 11770 78 11845 90
rect 11770 26 11781 78
rect 11833 26 11845 78
rect 11770 15 11845 26
rect 11675 -47 11750 -35
rect 11675 -99 11686 -47
rect 11738 -99 11750 -47
rect 11675 -110 11750 -99
rect 11780 -110 11830 15
rect 11925 -140 11975 120
rect 12150 78 12225 90
rect 12150 26 12161 78
rect 12213 26 12225 78
rect 12150 15 12225 26
rect 12164 -110 12215 15
rect 12255 -35 12306 90
rect 12340 78 12415 90
rect 12340 26 12351 78
rect 12403 26 12415 78
rect 12340 15 12415 26
rect 12245 -47 12320 -35
rect 12245 -99 12256 -47
rect 12308 -99 12320 -47
rect 12245 -110 12320 -99
rect 12350 -110 12402 15
rect 12450 -35 12501 90
rect 12535 78 12610 90
rect 12535 26 12546 78
rect 12598 26 12610 78
rect 12535 15 12610 26
rect 12435 -47 12510 -35
rect 12435 -99 12446 -47
rect 12498 -99 12510 -47
rect 12435 -110 12510 -99
rect 12545 -110 12596 15
rect 12685 -140 12740 120
rect 9900 -190 11975 -140
rect 12190 -190 12740 -140
rect 10205 -565 10600 -550
rect 10205 -1065 10216 -565
rect 10588 -1065 10600 -565
rect 10205 -1080 10600 -1065
rect 11925 -1260 11975 -190
rect 12200 -195 12740 -190
rect 12140 -558 12570 -525
rect 12140 -1058 12169 -558
rect 12541 -1058 12570 -558
rect 12140 -1090 12570 -1058
rect 12900 -1255 12955 120
rect 13365 -1260 13415 470
rect 15855 465 21775 515
rect 15855 175 15905 465
rect 13535 120 15625 170
rect 15855 125 21775 175
rect 13535 -145 13585 120
rect 13690 78 13765 90
rect 13690 26 13701 78
rect 13753 26 13765 78
rect 13690 15 13765 26
rect 13704 -30 13750 15
rect 13704 -98 13710 -30
rect 13744 -98 13750 -30
rect 13800 -35 13846 90
rect 13880 78 13955 90
rect 13880 26 13891 78
rect 13943 26 13955 78
rect 13880 15 13955 26
rect 13704 -110 13750 -98
rect 13785 -47 13860 -35
rect 13785 -99 13796 -47
rect 13848 -99 13860 -47
rect 13785 -110 13860 -99
rect 13895 -110 13942 15
rect 13990 -35 14038 90
rect 14075 78 14150 90
rect 14075 26 14086 78
rect 14138 26 14150 78
rect 14075 15 14150 26
rect 13975 -47 14050 -35
rect 13975 -99 13986 -47
rect 14038 -99 14050 -47
rect 13975 -110 14050 -99
rect 14085 -110 14134 15
rect 14184 -35 14231 90
rect 14265 78 14340 90
rect 14265 26 14276 78
rect 14328 26 14340 78
rect 14265 15 14340 26
rect 14170 -47 14245 -35
rect 14170 -99 14181 -47
rect 14233 -99 14245 -47
rect 14170 -110 14245 -99
rect 14280 -110 14326 15
rect 14375 -35 14422 90
rect 14460 78 14535 90
rect 14460 26 14471 78
rect 14523 26 14535 78
rect 14460 15 14535 26
rect 14360 -47 14435 -35
rect 14360 -99 14371 -47
rect 14423 -99 14435 -47
rect 14360 -110 14435 -99
rect 14470 -110 14518 15
rect 14565 -35 14614 90
rect 14645 78 14720 90
rect 14645 26 14656 78
rect 14708 26 14720 78
rect 14645 15 14720 26
rect 14550 -47 14625 -35
rect 14550 -99 14561 -47
rect 14613 -99 14625 -47
rect 14550 -110 14625 -99
rect 14664 -110 14711 15
rect 14760 -35 14806 90
rect 14840 78 14915 90
rect 14840 26 14851 78
rect 14903 26 14915 78
rect 14840 15 14915 26
rect 14745 -47 14820 -35
rect 14745 -99 14756 -47
rect 14808 -99 14820 -47
rect 14745 -110 14820 -99
rect 14855 -110 14902 15
rect 14950 -35 14998 90
rect 15030 78 15105 90
rect 15030 26 15041 78
rect 15093 26 15105 78
rect 15030 15 15105 26
rect 14935 -47 15010 -35
rect 14935 -99 14946 -47
rect 14998 -99 15010 -47
rect 14935 -110 15010 -99
rect 15048 -110 15096 15
rect 15144 -35 15191 90
rect 15225 78 15300 90
rect 15225 26 15236 78
rect 15288 26 15300 78
rect 15225 15 15300 26
rect 15130 -47 15205 -35
rect 15130 -99 15141 -47
rect 15193 -99 15205 -47
rect 15130 -110 15205 -99
rect 15240 -110 15286 15
rect 15335 -35 15382 90
rect 15415 78 15490 90
rect 15415 26 15426 78
rect 15478 26 15490 78
rect 15415 15 15490 26
rect 15320 -47 15395 -35
rect 15320 -99 15331 -47
rect 15383 -99 15395 -47
rect 15320 -110 15395 -99
rect 15430 -110 15478 15
rect 15525 -35 15574 90
rect 15610 78 15685 90
rect 15610 26 15621 78
rect 15673 26 15685 78
rect 15610 15 15685 26
rect 15510 -47 15585 -35
rect 15510 -99 15521 -47
rect 15573 -99 15585 -47
rect 15510 -110 15585 -99
rect 15624 -110 15671 15
rect 15855 -140 15905 125
rect 16046 122 16104 125
rect 16238 122 16296 125
rect 16430 122 16488 125
rect 16622 122 16680 125
rect 16814 122 16872 125
rect 17006 122 17064 125
rect 17198 122 17256 125
rect 17390 122 17448 125
rect 17582 122 17640 125
rect 17774 122 17832 125
rect 17966 122 18024 125
rect 18158 122 18216 125
rect 18350 122 18408 125
rect 18542 122 18600 125
rect 18734 122 18792 125
rect 18926 122 18984 125
rect 19118 122 19176 125
rect 19310 122 19368 125
rect 19502 122 19560 125
rect 19694 122 19752 125
rect 19886 122 19944 125
rect 20078 122 20136 125
rect 20270 122 20328 125
rect 20462 122 20520 125
rect 20654 122 20712 125
rect 20846 122 20904 125
rect 21038 122 21096 125
rect 21230 122 21288 125
rect 21422 122 21480 125
rect 21614 122 21672 125
rect 15985 78 16060 90
rect 15985 26 15996 78
rect 16048 26 16060 78
rect 15985 15 16060 26
rect 16004 -110 16050 15
rect 16100 -35 16146 90
rect 16175 78 16250 90
rect 16175 26 16186 78
rect 16238 26 16250 78
rect 16175 15 16250 26
rect 16085 -47 16160 -35
rect 16085 -99 16096 -47
rect 16148 -99 16160 -47
rect 16085 -110 16160 -99
rect 16195 -110 16242 15
rect 16290 -35 16338 90
rect 16370 78 16445 90
rect 16370 26 16381 78
rect 16433 26 16445 78
rect 16370 15 16445 26
rect 16275 -47 16350 -35
rect 16275 -99 16286 -47
rect 16338 -99 16350 -47
rect 16275 -110 16350 -99
rect 16385 -110 16434 15
rect 16484 -35 16530 90
rect 16565 78 16640 90
rect 16565 26 16576 78
rect 16628 26 16640 78
rect 16565 15 16640 26
rect 16470 -47 16545 -35
rect 16470 -99 16481 -47
rect 16533 -99 16545 -47
rect 16470 -110 16545 -99
rect 16580 -110 16626 15
rect 16675 -35 16722 90
rect 16755 78 16830 90
rect 16755 26 16766 78
rect 16818 26 16830 78
rect 16755 15 16830 26
rect 16660 -47 16735 -35
rect 16660 -99 16671 -47
rect 16723 -99 16735 -47
rect 16660 -110 16735 -99
rect 16770 -110 16818 15
rect 16868 -35 16915 90
rect 16950 78 17025 90
rect 16950 26 16961 78
rect 17013 26 17025 78
rect 16950 15 17025 26
rect 16855 -47 16930 -35
rect 16855 -99 16866 -47
rect 16918 -99 16930 -47
rect 16855 -110 16930 -99
rect 16964 -110 17010 15
rect 17060 -35 17106 90
rect 17140 78 17215 90
rect 17140 26 17151 78
rect 17203 26 17215 78
rect 17140 15 17215 26
rect 17040 -47 17115 -35
rect 17040 -99 17051 -47
rect 17103 -99 17115 -47
rect 17040 -110 17115 -99
rect 17155 -110 17202 15
rect 17250 -35 17298 90
rect 17335 78 17410 90
rect 17335 26 17346 78
rect 17398 26 17410 78
rect 17335 15 17410 26
rect 17240 -47 17315 -35
rect 17240 -99 17251 -47
rect 17303 -99 17315 -47
rect 17240 -110 17315 -99
rect 17348 -110 17395 15
rect 17444 -35 17490 90
rect 17525 78 17600 90
rect 17525 26 17536 78
rect 17588 26 17600 78
rect 17525 15 17600 26
rect 17425 -47 17500 -35
rect 17425 -99 17436 -47
rect 17488 -99 17500 -47
rect 17425 -110 17500 -99
rect 17540 -110 17586 15
rect 17635 -35 17682 90
rect 17715 78 17790 90
rect 17715 26 17726 78
rect 17778 26 17790 78
rect 17715 15 17790 26
rect 17620 -47 17695 -35
rect 17620 -99 17631 -47
rect 17683 -99 17695 -47
rect 17620 -110 17695 -99
rect 17732 -110 17780 15
rect 17828 -35 17875 90
rect 17910 78 17985 90
rect 17910 26 17921 78
rect 17973 26 17985 78
rect 17910 15 17985 26
rect 17815 -47 17890 -35
rect 17815 -99 17826 -47
rect 17878 -99 17890 -47
rect 17815 -110 17890 -99
rect 17924 -110 17970 15
rect 18020 -35 18066 90
rect 18100 78 18175 90
rect 18100 26 18111 78
rect 18163 26 18175 78
rect 18100 15 18175 26
rect 18000 -47 18075 -35
rect 18000 -99 18011 -47
rect 18063 -99 18075 -47
rect 18000 -110 18075 -99
rect 18115 -110 18162 15
rect 18210 -35 18258 90
rect 18295 78 18370 90
rect 18295 26 18306 78
rect 18358 26 18370 78
rect 18295 15 18370 26
rect 18195 -47 18270 -35
rect 18195 -99 18206 -47
rect 18258 -99 18270 -47
rect 18195 -110 18270 -99
rect 18308 -110 18355 15
rect 18404 -35 18450 90
rect 18485 78 18560 90
rect 18485 26 18496 78
rect 18548 26 18560 78
rect 18485 15 18560 26
rect 18385 -47 18460 -35
rect 18385 -99 18396 -47
rect 18448 -99 18460 -47
rect 18385 -110 18460 -99
rect 18500 -110 18546 15
rect 18595 -35 18642 90
rect 18675 78 18750 90
rect 18675 26 18686 78
rect 18738 26 18750 78
rect 18675 15 18750 26
rect 18580 -47 18655 -35
rect 18580 -99 18591 -47
rect 18643 -99 18655 -47
rect 18580 -110 18655 -99
rect 18690 -110 18738 15
rect 18788 -35 18835 90
rect 18870 78 18945 90
rect 18870 26 18881 78
rect 18933 26 18945 78
rect 18870 15 18945 26
rect 18770 -47 18845 -35
rect 18770 -99 18781 -47
rect 18833 -99 18845 -47
rect 18770 -110 18845 -99
rect 18884 -110 18930 15
rect 18980 -35 19026 90
rect 19060 78 19135 90
rect 19060 26 19071 78
rect 19123 26 19135 78
rect 19060 15 19135 26
rect 18965 -47 19040 -35
rect 18965 -99 18976 -47
rect 19028 -99 19040 -47
rect 18965 -110 19040 -99
rect 19075 -110 19122 15
rect 19170 -35 19218 90
rect 19255 78 19330 90
rect 19255 26 19266 78
rect 19318 26 19330 78
rect 19255 15 19330 26
rect 19155 -47 19230 -35
rect 19155 -99 19166 -47
rect 19218 -99 19230 -47
rect 19155 -110 19230 -99
rect 19268 -110 19315 15
rect 19364 -35 19410 90
rect 19445 78 19520 90
rect 19445 26 19456 78
rect 19508 26 19520 78
rect 19445 15 19520 26
rect 19350 -47 19425 -35
rect 19350 -99 19361 -47
rect 19413 -99 19425 -47
rect 19350 -110 19425 -99
rect 19460 -110 19506 15
rect 19555 -35 19602 90
rect 19635 78 19710 90
rect 19635 26 19646 78
rect 19698 26 19710 78
rect 19635 15 19710 26
rect 19540 -47 19615 -35
rect 19540 -99 19551 -47
rect 19603 -99 19615 -47
rect 19540 -110 19615 -99
rect 19650 -110 19698 15
rect 19748 -35 19795 90
rect 19830 78 19905 90
rect 19830 26 19841 78
rect 19893 26 19905 78
rect 19830 15 19905 26
rect 19735 -47 19810 -35
rect 19735 -99 19746 -47
rect 19798 -99 19810 -47
rect 19735 -110 19810 -99
rect 19844 -110 19890 15
rect 19940 -35 19986 90
rect 20020 78 20095 90
rect 20020 26 20031 78
rect 20083 26 20095 78
rect 20020 15 20095 26
rect 19925 -47 20000 -35
rect 19925 -99 19936 -47
rect 19988 -99 20000 -47
rect 19925 -110 20000 -99
rect 20035 -110 20082 15
rect 20132 -35 20180 90
rect 20215 78 20290 90
rect 20215 26 20226 78
rect 20278 26 20290 78
rect 20215 15 20290 26
rect 20115 -47 20190 -35
rect 20115 -99 20126 -47
rect 20178 -99 20190 -47
rect 20115 -110 20190 -99
rect 20228 -110 20275 15
rect 20324 -35 20370 90
rect 20405 78 20480 90
rect 20405 26 20416 78
rect 20468 26 20480 78
rect 20405 15 20480 26
rect 20310 -47 20385 -35
rect 20310 -99 20321 -47
rect 20373 -99 20385 -47
rect 20310 -110 20385 -99
rect 20420 -110 20466 15
rect 20515 -35 20562 90
rect 20600 78 20675 90
rect 20600 26 20611 78
rect 20663 26 20675 78
rect 20600 15 20675 26
rect 20500 -47 20575 -35
rect 20500 -99 20511 -47
rect 20563 -99 20575 -47
rect 20500 -110 20575 -99
rect 20610 -110 20658 15
rect 20708 -35 20755 90
rect 20790 78 20865 90
rect 20790 26 20801 78
rect 20853 26 20865 78
rect 20790 15 20865 26
rect 20695 -47 20770 -35
rect 20695 -99 20706 -47
rect 20758 -99 20770 -47
rect 20695 -110 20770 -99
rect 20804 -110 20850 15
rect 20900 -35 20946 90
rect 20980 78 21055 90
rect 20980 26 20991 78
rect 21043 26 21055 78
rect 20980 15 21055 26
rect 20885 -47 20960 -35
rect 20885 -99 20896 -47
rect 20948 -99 20960 -47
rect 20885 -110 20960 -99
rect 20995 -110 21042 15
rect 21090 -35 21138 90
rect 21175 78 21250 90
rect 21175 26 21186 78
rect 21238 26 21250 78
rect 21175 15 21250 26
rect 21075 -47 21150 -35
rect 21075 -99 21086 -47
rect 21138 -99 21150 -47
rect 21075 -110 21150 -99
rect 21188 -110 21235 15
rect 21284 -35 21330 90
rect 21365 78 21440 90
rect 21365 26 21376 78
rect 21428 26 21440 78
rect 21365 15 21440 26
rect 21270 -47 21345 -35
rect 21270 -99 21281 -47
rect 21333 -99 21345 -47
rect 21270 -110 21345 -99
rect 21380 -110 21426 15
rect 21475 -35 21522 90
rect 21555 78 21630 90
rect 21555 26 21566 78
rect 21618 26 21630 78
rect 21555 15 21630 26
rect 21460 -47 21535 -35
rect 21460 -99 21471 -47
rect 21523 -99 21535 -47
rect 21460 -110 21535 -99
rect 21570 -110 21618 15
rect 21668 -35 21715 90
rect 21750 78 21825 90
rect 21750 26 21761 78
rect 21813 26 21825 78
rect 21750 15 21825 26
rect 21650 -47 21725 -35
rect 21650 -99 21661 -47
rect 21713 -99 21725 -47
rect 21650 -110 21725 -99
rect 21764 -110 21810 15
rect 13842 -145 13900 -142
rect 14034 -145 14092 -142
rect 14226 -145 14284 -142
rect 14418 -145 14476 -142
rect 14610 -145 14668 -142
rect 14802 -145 14860 -142
rect 14994 -145 15052 -142
rect 15186 -145 15244 -142
rect 15378 -145 15436 -142
rect 15570 -145 15628 -142
rect 13515 -157 15675 -145
rect 13515 -209 13526 -157
rect 13578 -195 15675 -157
rect 15855 -190 21775 -140
rect 13578 -209 13590 -195
rect 13515 -220 13590 -209
rect 13750 -570 14135 -560
rect 13750 -1646 13756 -570
rect 14128 -1646 14135 -570
rect 13750 -1655 14135 -1646
rect 15855 -1840 15905 -190
rect 17435 -572 17870 -530
rect 17435 -1648 17466 -572
rect 17838 -1648 17870 -572
rect 17435 -1675 17870 -1648
<< via1 >>
rect 10221 1205 10593 1705
rect 12186 1202 12558 1702
rect 13744 1197 14116 2273
rect 17461 1197 17833 2273
rect 13526 796 13578 848
rect 9956 686 10008 738
rect 9861 561 9913 613
rect 10151 686 10203 738
rect 10051 561 10103 613
rect 10341 686 10393 738
rect 10241 561 10293 613
rect 10531 686 10583 738
rect 10431 561 10483 613
rect 10721 686 10773 738
rect 10631 561 10683 613
rect 10911 686 10963 738
rect 10821 561 10873 613
rect 11106 686 11158 738
rect 11016 561 11068 613
rect 11301 686 11353 738
rect 11206 561 11258 613
rect 11491 686 11543 738
rect 11396 561 11448 613
rect 11686 686 11738 738
rect 11591 561 11643 613
rect 11781 561 11833 613
rect 12256 686 12308 738
rect 12161 561 12213 613
rect 12446 686 12498 738
rect 12351 561 12403 613
rect 12546 561 12598 613
rect 13796 686 13848 738
rect 13701 561 13753 613
rect 13986 686 14038 738
rect 13891 561 13943 613
rect 14181 686 14233 738
rect 14086 561 14138 613
rect 14371 686 14423 738
rect 14276 561 14328 613
rect 14561 686 14613 738
rect 14471 561 14523 613
rect 14756 686 14808 738
rect 14656 561 14708 613
rect 14946 686 14998 738
rect 14851 561 14903 613
rect 15141 686 15193 738
rect 15041 561 15093 613
rect 15331 686 15383 738
rect 15236 561 15288 613
rect 15521 686 15573 738
rect 15426 561 15478 613
rect 15621 561 15673 613
rect 16096 686 16148 738
rect 15996 561 16048 613
rect 16286 686 16338 738
rect 16186 561 16238 613
rect 16481 686 16533 738
rect 16381 561 16433 613
rect 16671 686 16723 738
rect 16576 561 16628 613
rect 16866 686 16918 738
rect 16766 561 16818 613
rect 17051 686 17103 738
rect 16961 561 17013 613
rect 17251 686 17303 738
rect 17151 561 17203 613
rect 17436 686 17488 738
rect 17346 561 17398 613
rect 17631 686 17683 738
rect 17536 561 17588 613
rect 17826 686 17878 738
rect 17726 561 17778 613
rect 18011 686 18063 738
rect 17921 561 17973 613
rect 18206 686 18258 738
rect 18111 561 18163 613
rect 18396 686 18448 738
rect 18306 561 18358 613
rect 18591 686 18643 738
rect 18496 561 18548 613
rect 18781 686 18833 738
rect 18686 561 18738 613
rect 18976 686 19028 738
rect 18881 561 18933 613
rect 19166 686 19218 738
rect 19071 561 19123 613
rect 19361 686 19413 738
rect 19266 561 19318 613
rect 19551 686 19603 738
rect 19456 561 19508 613
rect 19746 686 19798 738
rect 19646 561 19698 613
rect 19936 686 19988 738
rect 19841 561 19893 613
rect 20126 686 20178 738
rect 20031 561 20083 613
rect 20321 686 20373 738
rect 20226 561 20278 613
rect 20511 686 20563 738
rect 20416 561 20468 613
rect 20706 686 20758 738
rect 20611 561 20663 613
rect 20896 686 20948 738
rect 20801 561 20853 613
rect 21086 686 21138 738
rect 20991 561 21043 613
rect 21281 686 21333 738
rect 21186 561 21238 613
rect 21471 686 21523 738
rect 21376 561 21428 613
rect 21661 686 21713 738
rect 21566 561 21618 613
rect 21761 561 21813 613
rect 9861 26 9913 78
rect 10051 26 10103 78
rect 9956 -99 10008 -47
rect 10241 26 10293 78
rect 10151 -99 10203 -47
rect 10431 26 10483 78
rect 10341 -99 10393 -47
rect 10631 26 10683 78
rect 10531 -99 10583 -47
rect 10821 26 10873 78
rect 10721 -99 10773 -47
rect 11016 26 11068 78
rect 10911 -99 10963 -47
rect 11206 26 11258 78
rect 11106 -99 11158 -47
rect 11396 26 11448 78
rect 11301 -99 11353 -47
rect 11591 26 11643 78
rect 11491 -99 11543 -47
rect 11781 26 11833 78
rect 11686 -99 11738 -47
rect 12161 26 12213 78
rect 12351 26 12403 78
rect 12256 -99 12308 -47
rect 12546 26 12598 78
rect 12446 -99 12498 -47
rect 10216 -1065 10588 -565
rect 12169 -1058 12541 -558
rect 13701 26 13753 78
rect 13891 26 13943 78
rect 13796 -99 13848 -47
rect 14086 26 14138 78
rect 13986 -99 14038 -47
rect 14276 26 14328 78
rect 14181 -99 14233 -47
rect 14471 26 14523 78
rect 14371 -99 14423 -47
rect 14656 26 14708 78
rect 14561 -99 14613 -47
rect 14851 26 14903 78
rect 14756 -99 14808 -47
rect 15041 26 15093 78
rect 14946 -99 14998 -47
rect 15236 26 15288 78
rect 15141 -99 15193 -47
rect 15426 26 15478 78
rect 15331 -99 15383 -47
rect 15621 26 15673 78
rect 15521 -99 15573 -47
rect 15996 26 16048 78
rect 16186 26 16238 78
rect 16096 -99 16148 -47
rect 16381 26 16433 78
rect 16286 -99 16338 -47
rect 16576 26 16628 78
rect 16481 -99 16533 -47
rect 16766 26 16818 78
rect 16671 -99 16723 -47
rect 16961 26 17013 78
rect 16866 -99 16918 -47
rect 17151 26 17203 78
rect 17051 -99 17103 -47
rect 17346 26 17398 78
rect 17251 -99 17303 -47
rect 17536 26 17588 78
rect 17436 -99 17488 -47
rect 17726 26 17778 78
rect 17631 -99 17683 -47
rect 17921 26 17973 78
rect 17826 -99 17878 -47
rect 18111 26 18163 78
rect 18011 -99 18063 -47
rect 18306 26 18358 78
rect 18206 -99 18258 -47
rect 18496 26 18548 78
rect 18396 -99 18448 -47
rect 18686 26 18738 78
rect 18591 -99 18643 -47
rect 18881 26 18933 78
rect 18781 -99 18833 -47
rect 19071 26 19123 78
rect 18976 -99 19028 -47
rect 19266 26 19318 78
rect 19166 -99 19218 -47
rect 19456 26 19508 78
rect 19361 -99 19413 -47
rect 19646 26 19698 78
rect 19551 -99 19603 -47
rect 19841 26 19893 78
rect 19746 -99 19798 -47
rect 20031 26 20083 78
rect 19936 -99 19988 -47
rect 20226 26 20278 78
rect 20126 -99 20178 -47
rect 20416 26 20468 78
rect 20321 -99 20373 -47
rect 20611 26 20663 78
rect 20511 -99 20563 -47
rect 20801 26 20853 78
rect 20706 -99 20758 -47
rect 20991 26 21043 78
rect 20896 -99 20948 -47
rect 21186 26 21238 78
rect 21086 -99 21138 -47
rect 21376 26 21428 78
rect 21281 -99 21333 -47
rect 21566 26 21618 78
rect 21471 -99 21523 -47
rect 21761 26 21813 78
rect 21661 -99 21713 -47
rect 13526 -209 13578 -157
rect 13756 -1646 14128 -570
rect 17466 -1648 17838 -572
<< metal2 >>
rect 13715 2273 14160 2315
rect 13715 2243 13744 2273
rect 14116 2243 14160 2273
rect 10195 1705 10620 1735
rect 10195 1683 10221 1705
rect 10593 1683 10620 1705
rect 10195 1227 10219 1683
rect 10595 1227 10620 1683
rect 10195 1205 10221 1227
rect 10593 1205 10620 1227
rect 10195 1165 10620 1205
rect 12155 1702 12590 1735
rect 12155 1202 12186 1702
rect 12558 1202 12590 1702
rect 12155 1070 12590 1202
rect 13715 1227 13742 2243
rect 14118 1227 14160 2243
rect 13715 1197 13744 1227
rect 14116 1197 14160 1227
rect 13715 1165 14160 1197
rect 17435 2273 17870 2310
rect 17435 2243 17461 2273
rect 17833 2243 17870 2273
rect 17435 1227 17459 2243
rect 17835 1227 17870 2243
rect 17435 1197 17461 1227
rect 17833 1197 17870 1227
rect 17435 1165 17870 1197
rect 12155 1000 13585 1070
rect 8845 975 9985 980
rect 8845 738 11835 975
rect 8845 686 9956 738
rect 10008 686 10151 738
rect 10203 686 10341 738
rect 10393 686 10531 738
rect 10583 686 10721 738
rect 10773 686 10911 738
rect 10963 686 11106 738
rect 11158 686 11301 738
rect 11353 686 11491 738
rect 11543 686 11686 738
rect 11738 686 11835 738
rect 8845 680 11835 686
rect 12155 738 12590 1000
rect 13515 860 13585 1000
rect 13515 848 13590 860
rect 13515 796 13526 848
rect 13578 796 13590 848
rect 13515 785 13590 796
rect 12155 686 12256 738
rect 12308 686 12446 738
rect 12498 686 12590 738
rect 8845 -40 9445 680
rect 12155 675 12590 686
rect 13785 758 13860 775
rect 13785 738 13797 758
rect 13785 686 13796 738
rect 13853 702 13860 758
rect 13848 686 13860 702
rect 13785 675 13860 686
rect 13975 758 14050 775
rect 13975 738 13987 758
rect 13975 686 13986 738
rect 14043 702 14050 758
rect 14038 686 14050 702
rect 13975 675 14050 686
rect 14170 758 14245 775
rect 14170 738 14182 758
rect 14170 686 14181 738
rect 14238 702 14245 758
rect 14233 686 14245 702
rect 14170 675 14245 686
rect 14360 758 14435 775
rect 14360 738 14372 758
rect 14360 686 14371 738
rect 14428 702 14435 758
rect 14423 686 14435 702
rect 14360 675 14435 686
rect 14550 758 14625 775
rect 14550 738 14562 758
rect 14550 686 14561 738
rect 14618 702 14625 758
rect 14613 686 14625 702
rect 14550 675 14625 686
rect 14745 758 14820 775
rect 14745 738 14757 758
rect 14745 686 14756 738
rect 14813 702 14820 758
rect 14808 686 14820 702
rect 14745 675 14820 686
rect 14935 758 15010 775
rect 14935 738 14947 758
rect 14935 686 14946 738
rect 15003 702 15010 758
rect 14998 686 15010 702
rect 14935 675 15010 686
rect 15130 758 15205 775
rect 15130 738 15142 758
rect 15130 686 15141 738
rect 15198 702 15205 758
rect 15193 686 15205 702
rect 15130 675 15205 686
rect 15320 758 15395 775
rect 15320 738 15332 758
rect 15320 686 15331 738
rect 15388 702 15395 758
rect 15383 686 15395 702
rect 15320 675 15395 686
rect 15510 758 15585 775
rect 15510 738 15522 758
rect 15510 686 15521 738
rect 15578 702 15585 758
rect 15573 686 15585 702
rect 15510 675 15585 686
rect 16085 758 16160 775
rect 16085 702 16092 758
rect 16085 686 16096 702
rect 16148 686 16160 758
rect 16085 675 16160 686
rect 16275 758 16350 775
rect 16275 702 16282 758
rect 16275 686 16286 702
rect 16338 686 16350 758
rect 16275 675 16350 686
rect 16470 758 16545 775
rect 16470 702 16477 758
rect 16470 686 16481 702
rect 16533 686 16545 758
rect 16470 675 16545 686
rect 16660 758 16735 775
rect 16660 702 16667 758
rect 16660 686 16671 702
rect 16723 686 16735 758
rect 16660 675 16735 686
rect 16855 758 16930 775
rect 16855 702 16862 758
rect 16855 686 16866 702
rect 16918 686 16930 758
rect 16855 675 16930 686
rect 17040 758 17115 775
rect 17040 702 17047 758
rect 17040 686 17051 702
rect 17103 686 17115 758
rect 17040 675 17115 686
rect 17240 758 17315 775
rect 17240 702 17247 758
rect 17240 686 17251 702
rect 17303 686 17315 758
rect 17240 675 17315 686
rect 17425 758 17500 775
rect 17425 702 17432 758
rect 17425 686 17436 702
rect 17488 686 17500 758
rect 17425 675 17500 686
rect 17620 758 17695 775
rect 17620 702 17627 758
rect 17620 686 17631 702
rect 17683 686 17695 758
rect 17620 675 17695 686
rect 17815 758 17890 775
rect 17815 702 17822 758
rect 17815 686 17826 702
rect 17878 686 17890 758
rect 17815 675 17890 686
rect 18000 758 18075 775
rect 18000 702 18007 758
rect 18000 686 18011 702
rect 18063 686 18075 758
rect 18000 675 18075 686
rect 18195 758 18270 775
rect 18195 702 18202 758
rect 18195 686 18206 702
rect 18258 686 18270 758
rect 18195 675 18270 686
rect 18385 758 18460 775
rect 18385 702 18392 758
rect 18385 686 18396 702
rect 18448 686 18460 758
rect 18385 675 18460 686
rect 18580 758 18655 775
rect 18580 702 18587 758
rect 18580 686 18591 702
rect 18643 686 18655 758
rect 18580 675 18655 686
rect 18770 758 18845 775
rect 18770 702 18777 758
rect 18770 686 18781 702
rect 18833 686 18845 758
rect 18770 675 18845 686
rect 18965 758 19040 775
rect 18965 702 18972 758
rect 18965 686 18976 702
rect 19028 686 19040 758
rect 18965 675 19040 686
rect 19155 758 19230 775
rect 19155 702 19162 758
rect 19155 686 19166 702
rect 19218 686 19230 758
rect 19155 675 19230 686
rect 19350 758 19425 775
rect 19350 702 19357 758
rect 19350 686 19361 702
rect 19413 686 19425 758
rect 19350 675 19425 686
rect 19540 758 19615 775
rect 19540 702 19547 758
rect 19540 686 19551 702
rect 19603 686 19615 758
rect 19540 675 19615 686
rect 19735 758 19810 775
rect 19735 702 19742 758
rect 19735 686 19746 702
rect 19798 686 19810 758
rect 19735 675 19810 686
rect 19925 758 20000 775
rect 19925 702 19932 758
rect 19925 686 19936 702
rect 19988 686 20000 758
rect 19925 675 20000 686
rect 20115 758 20190 775
rect 20115 702 20122 758
rect 20115 686 20126 702
rect 20178 686 20190 758
rect 20115 675 20190 686
rect 20310 758 20385 775
rect 20310 702 20317 758
rect 20310 686 20321 702
rect 20373 686 20385 758
rect 20310 675 20385 686
rect 20500 758 20575 775
rect 20500 702 20507 758
rect 20500 686 20511 702
rect 20563 686 20575 758
rect 20500 675 20575 686
rect 20695 758 20770 775
rect 20695 702 20702 758
rect 20695 686 20706 702
rect 20758 686 20770 758
rect 20695 675 20770 686
rect 20885 758 20960 775
rect 20885 702 20892 758
rect 20885 686 20896 702
rect 20948 686 20960 758
rect 20885 675 20960 686
rect 21075 758 21150 775
rect 21075 702 21082 758
rect 21075 686 21086 702
rect 21138 686 21150 758
rect 21075 675 21150 686
rect 21270 758 21345 775
rect 21270 702 21277 758
rect 21270 686 21281 702
rect 21333 686 21345 758
rect 21270 675 21345 686
rect 21460 758 21535 775
rect 21460 702 21467 758
rect 21460 686 21471 702
rect 21523 686 21535 758
rect 21460 675 21535 686
rect 21650 758 21725 775
rect 21650 702 21657 758
rect 21650 686 21661 702
rect 21713 686 21725 758
rect 21650 675 21725 686
rect 12150 620 12225 625
rect 12340 620 12415 625
rect 12535 620 12610 625
rect 9850 613 12610 620
rect 9850 561 9861 613
rect 9913 561 10051 613
rect 10103 561 10241 613
rect 10293 561 10431 613
rect 10483 561 10631 613
rect 10683 561 10821 613
rect 10873 561 11016 613
rect 11068 561 11206 613
rect 11258 561 11396 613
rect 11448 561 11591 613
rect 11643 561 11781 613
rect 11833 561 12161 613
rect 12213 561 12351 613
rect 12403 561 12546 613
rect 12598 561 12610 613
rect 9850 78 12610 561
rect 13690 613 13765 625
rect 13690 561 13701 613
rect 13753 598 13765 613
rect 13690 542 13702 561
rect 13758 542 13765 598
rect 13690 525 13765 542
rect 13880 613 13955 625
rect 13880 561 13891 613
rect 13943 598 13955 613
rect 13880 542 13892 561
rect 13948 542 13955 598
rect 13880 525 13955 542
rect 14075 613 14150 625
rect 14075 561 14086 613
rect 14138 598 14150 613
rect 14075 542 14087 561
rect 14143 542 14150 598
rect 14075 525 14150 542
rect 14265 613 14340 625
rect 14265 561 14276 613
rect 14328 598 14340 613
rect 14265 542 14277 561
rect 14333 542 14340 598
rect 14265 525 14340 542
rect 14460 613 14535 625
rect 14460 561 14471 613
rect 14523 598 14535 613
rect 14460 542 14472 561
rect 14528 542 14535 598
rect 14460 525 14535 542
rect 14645 613 14720 625
rect 14645 561 14656 613
rect 14708 598 14720 613
rect 14645 542 14657 561
rect 14713 542 14720 598
rect 14645 525 14720 542
rect 14840 613 14915 625
rect 14840 561 14851 613
rect 14903 598 14915 613
rect 14840 542 14852 561
rect 14908 542 14915 598
rect 14840 525 14915 542
rect 15030 613 15105 625
rect 15030 561 15041 613
rect 15093 598 15105 613
rect 15030 542 15042 561
rect 15098 542 15105 598
rect 15030 525 15105 542
rect 15225 613 15300 625
rect 15225 561 15236 613
rect 15288 598 15300 613
rect 15225 542 15237 561
rect 15293 542 15300 598
rect 15225 525 15300 542
rect 15415 613 15490 625
rect 15415 561 15426 613
rect 15478 598 15490 613
rect 15415 542 15427 561
rect 15483 542 15490 598
rect 15415 525 15490 542
rect 15610 613 15685 625
rect 15610 561 15621 613
rect 15673 598 15685 613
rect 15610 542 15622 561
rect 15678 542 15685 598
rect 15610 525 15685 542
rect 15985 613 16060 625
rect 15985 561 15996 613
rect 16048 598 16060 613
rect 15985 542 15997 561
rect 16053 542 16060 598
rect 15985 525 16060 542
rect 16175 613 16250 625
rect 16175 561 16186 613
rect 16238 598 16250 613
rect 16175 542 16187 561
rect 16243 542 16250 598
rect 16175 525 16250 542
rect 16370 613 16445 625
rect 16370 561 16381 613
rect 16433 598 16445 613
rect 16370 542 16382 561
rect 16438 542 16445 598
rect 16370 525 16445 542
rect 16565 613 16640 625
rect 16565 561 16576 613
rect 16628 598 16640 613
rect 16565 542 16577 561
rect 16633 542 16640 598
rect 16565 525 16640 542
rect 16755 613 16830 625
rect 16755 561 16766 613
rect 16818 598 16830 613
rect 16755 542 16767 561
rect 16823 542 16830 598
rect 16755 525 16830 542
rect 16950 613 17025 625
rect 16950 561 16961 613
rect 17013 598 17025 613
rect 16950 542 16962 561
rect 17018 542 17025 598
rect 16950 525 17025 542
rect 17140 613 17215 625
rect 17140 561 17151 613
rect 17203 598 17215 613
rect 17140 542 17152 561
rect 17208 542 17215 598
rect 17140 525 17215 542
rect 17335 613 17410 625
rect 17335 561 17346 613
rect 17398 598 17410 613
rect 17335 542 17347 561
rect 17403 542 17410 598
rect 17335 525 17410 542
rect 17525 613 17600 625
rect 17525 561 17536 613
rect 17588 598 17600 613
rect 17525 542 17537 561
rect 17593 542 17600 598
rect 17525 525 17600 542
rect 17715 613 17790 625
rect 17715 561 17726 613
rect 17778 598 17790 613
rect 17715 542 17727 561
rect 17783 542 17790 598
rect 17715 525 17790 542
rect 17910 613 17985 625
rect 17910 561 17921 613
rect 17973 598 17985 613
rect 17910 542 17922 561
rect 17978 542 17985 598
rect 17910 525 17985 542
rect 18100 613 18175 625
rect 18100 561 18111 613
rect 18163 598 18175 613
rect 18100 542 18112 561
rect 18168 542 18175 598
rect 18100 525 18175 542
rect 18295 613 18370 625
rect 18295 561 18306 613
rect 18358 598 18370 613
rect 18295 542 18307 561
rect 18363 542 18370 598
rect 18295 525 18370 542
rect 18485 613 18560 625
rect 18485 561 18496 613
rect 18548 598 18560 613
rect 18485 542 18497 561
rect 18553 542 18560 598
rect 18485 525 18560 542
rect 18675 613 18750 625
rect 18675 561 18686 613
rect 18738 598 18750 613
rect 18675 542 18687 561
rect 18743 542 18750 598
rect 18675 525 18750 542
rect 18870 613 18945 625
rect 18870 561 18881 613
rect 18933 598 18945 613
rect 18870 542 18882 561
rect 18938 542 18945 598
rect 18870 525 18945 542
rect 19060 613 19135 625
rect 19060 561 19071 613
rect 19123 598 19135 613
rect 19060 542 19072 561
rect 19128 542 19135 598
rect 19060 525 19135 542
rect 19255 613 19330 625
rect 19255 561 19266 613
rect 19318 598 19330 613
rect 19255 542 19267 561
rect 19323 542 19330 598
rect 19255 525 19330 542
rect 19445 613 19520 625
rect 19445 561 19456 613
rect 19508 598 19520 613
rect 19445 542 19457 561
rect 19513 542 19520 598
rect 19445 525 19520 542
rect 19635 613 19710 625
rect 19635 561 19646 613
rect 19698 598 19710 613
rect 19635 542 19647 561
rect 19703 542 19710 598
rect 19635 525 19710 542
rect 19830 613 19905 625
rect 19830 561 19841 613
rect 19893 598 19905 613
rect 19830 542 19842 561
rect 19898 542 19905 598
rect 19830 525 19905 542
rect 20020 613 20095 625
rect 20020 561 20031 613
rect 20083 598 20095 613
rect 20020 542 20032 561
rect 20088 542 20095 598
rect 20020 525 20095 542
rect 20215 613 20290 625
rect 20215 561 20226 613
rect 20278 598 20290 613
rect 20215 542 20227 561
rect 20283 542 20290 598
rect 20215 525 20290 542
rect 20405 613 20480 625
rect 20405 561 20416 613
rect 20468 598 20480 613
rect 20405 542 20417 561
rect 20473 542 20480 598
rect 20405 525 20480 542
rect 20600 613 20675 625
rect 20600 561 20611 613
rect 20663 598 20675 613
rect 20600 542 20612 561
rect 20668 542 20675 598
rect 20600 525 20675 542
rect 20790 613 20865 625
rect 20790 561 20801 613
rect 20853 598 20865 613
rect 20790 542 20802 561
rect 20858 542 20865 598
rect 20790 525 20865 542
rect 20980 613 21055 625
rect 20980 561 20991 613
rect 21043 598 21055 613
rect 20980 542 20992 561
rect 21048 542 21055 598
rect 20980 525 21055 542
rect 21175 613 21250 625
rect 21175 561 21186 613
rect 21238 598 21250 613
rect 21175 542 21187 561
rect 21243 542 21250 598
rect 21175 525 21250 542
rect 21365 613 21440 625
rect 21365 561 21376 613
rect 21428 598 21440 613
rect 21365 542 21377 561
rect 21433 542 21440 598
rect 21365 525 21440 542
rect 21555 613 21630 625
rect 21555 561 21566 613
rect 21618 598 21630 613
rect 21555 542 21567 561
rect 21623 542 21630 598
rect 21555 525 21630 542
rect 21750 613 21825 625
rect 21750 561 21761 613
rect 21813 598 21825 613
rect 21750 542 21762 561
rect 21818 542 21825 598
rect 21750 525 21825 542
rect 9850 26 9861 78
rect 9913 26 10051 78
rect 10103 26 10241 78
rect 10293 26 10431 78
rect 10483 26 10631 78
rect 10683 26 10821 78
rect 10873 26 11016 78
rect 11068 26 11206 78
rect 11258 26 11396 78
rect 11448 26 11591 78
rect 11643 26 11781 78
rect 11833 26 12161 78
rect 12213 26 12351 78
rect 12403 26 12546 78
rect 12598 26 12610 78
rect 9850 20 12610 26
rect 12150 15 12225 20
rect 12340 15 12415 20
rect 12535 15 12610 20
rect 13690 98 13765 115
rect 13690 78 13702 98
rect 13690 26 13701 78
rect 13758 42 13765 98
rect 13753 26 13765 42
rect 13690 15 13765 26
rect 13880 98 13955 115
rect 13880 78 13892 98
rect 13880 26 13891 78
rect 13948 42 13955 98
rect 13943 26 13955 42
rect 13880 15 13955 26
rect 14075 98 14150 115
rect 14075 78 14087 98
rect 14075 26 14086 78
rect 14143 42 14150 98
rect 14138 26 14150 42
rect 14075 15 14150 26
rect 14265 98 14340 115
rect 14265 78 14277 98
rect 14265 26 14276 78
rect 14333 42 14340 98
rect 14328 26 14340 42
rect 14265 15 14340 26
rect 14460 98 14535 115
rect 14460 78 14472 98
rect 14460 26 14471 78
rect 14528 42 14535 98
rect 14523 26 14535 42
rect 14460 15 14535 26
rect 14645 98 14720 115
rect 14645 78 14657 98
rect 14645 26 14656 78
rect 14713 42 14720 98
rect 14708 26 14720 42
rect 14645 15 14720 26
rect 14840 98 14915 115
rect 14840 78 14852 98
rect 14840 26 14851 78
rect 14908 42 14915 98
rect 14903 26 14915 42
rect 14840 15 14915 26
rect 15030 98 15105 115
rect 15030 78 15042 98
rect 15030 26 15041 78
rect 15098 42 15105 98
rect 15093 26 15105 42
rect 15030 15 15105 26
rect 15225 98 15300 115
rect 15225 78 15237 98
rect 15225 26 15236 78
rect 15293 42 15300 98
rect 15288 26 15300 42
rect 15225 15 15300 26
rect 15415 98 15490 115
rect 15415 78 15427 98
rect 15415 26 15426 78
rect 15483 42 15490 98
rect 15478 26 15490 42
rect 15415 15 15490 26
rect 15610 98 15685 115
rect 15610 78 15622 98
rect 15610 26 15621 78
rect 15678 42 15685 98
rect 15673 26 15685 42
rect 15610 15 15685 26
rect 15985 98 16060 115
rect 15985 78 15997 98
rect 15985 26 15996 78
rect 16053 42 16060 98
rect 16048 26 16060 42
rect 15985 15 16060 26
rect 16175 98 16250 115
rect 16175 78 16187 98
rect 16175 26 16186 78
rect 16243 42 16250 98
rect 16238 26 16250 42
rect 16175 15 16250 26
rect 16370 98 16445 115
rect 16370 78 16382 98
rect 16370 26 16381 78
rect 16438 42 16445 98
rect 16433 26 16445 42
rect 16370 15 16445 26
rect 16565 98 16640 115
rect 16565 78 16577 98
rect 16565 26 16576 78
rect 16633 42 16640 98
rect 16628 26 16640 42
rect 16565 15 16640 26
rect 16755 98 16830 115
rect 16755 78 16767 98
rect 16755 26 16766 78
rect 16823 42 16830 98
rect 16818 26 16830 42
rect 16755 15 16830 26
rect 16950 98 17025 115
rect 16950 78 16962 98
rect 16950 26 16961 78
rect 17018 42 17025 98
rect 17013 26 17025 42
rect 16950 15 17025 26
rect 17140 98 17215 115
rect 17140 78 17152 98
rect 17140 26 17151 78
rect 17208 42 17215 98
rect 17203 26 17215 42
rect 17140 15 17215 26
rect 17335 98 17410 115
rect 17335 78 17347 98
rect 17335 26 17346 78
rect 17403 42 17410 98
rect 17398 26 17410 42
rect 17335 15 17410 26
rect 17525 98 17600 115
rect 17525 78 17537 98
rect 17525 26 17536 78
rect 17593 42 17600 98
rect 17588 26 17600 42
rect 17525 15 17600 26
rect 17715 98 17790 115
rect 17715 78 17727 98
rect 17715 26 17726 78
rect 17783 42 17790 98
rect 17778 26 17790 42
rect 17715 15 17790 26
rect 17910 98 17985 115
rect 17910 78 17922 98
rect 17910 26 17921 78
rect 17978 42 17985 98
rect 17973 26 17985 42
rect 17910 15 17985 26
rect 18100 98 18175 115
rect 18100 78 18112 98
rect 18100 26 18111 78
rect 18168 42 18175 98
rect 18163 26 18175 42
rect 18100 15 18175 26
rect 18295 98 18370 115
rect 18295 78 18307 98
rect 18295 26 18306 78
rect 18363 42 18370 98
rect 18358 26 18370 42
rect 18295 15 18370 26
rect 18485 98 18560 115
rect 18485 78 18497 98
rect 18485 26 18496 78
rect 18553 42 18560 98
rect 18548 26 18560 42
rect 18485 15 18560 26
rect 18675 98 18750 115
rect 18675 78 18687 98
rect 18675 26 18686 78
rect 18743 42 18750 98
rect 18738 26 18750 42
rect 18675 15 18750 26
rect 18870 98 18945 115
rect 18870 78 18882 98
rect 18870 26 18881 78
rect 18938 42 18945 98
rect 18933 26 18945 42
rect 18870 15 18945 26
rect 19060 98 19135 115
rect 19060 78 19072 98
rect 19060 26 19071 78
rect 19128 42 19135 98
rect 19123 26 19135 42
rect 19060 15 19135 26
rect 19255 98 19330 115
rect 19255 78 19267 98
rect 19255 26 19266 78
rect 19323 42 19330 98
rect 19318 26 19330 42
rect 19255 15 19330 26
rect 19445 98 19520 115
rect 19445 78 19457 98
rect 19445 26 19456 78
rect 19513 42 19520 98
rect 19508 26 19520 42
rect 19445 15 19520 26
rect 19635 98 19710 115
rect 19635 78 19647 98
rect 19635 26 19646 78
rect 19703 42 19710 98
rect 19698 26 19710 42
rect 19635 15 19710 26
rect 19830 98 19905 115
rect 19830 78 19842 98
rect 19830 26 19841 78
rect 19898 42 19905 98
rect 19893 26 19905 42
rect 19830 15 19905 26
rect 20020 98 20095 115
rect 20020 78 20032 98
rect 20020 26 20031 78
rect 20088 42 20095 98
rect 20083 26 20095 42
rect 20020 15 20095 26
rect 20215 98 20290 115
rect 20215 78 20227 98
rect 20215 26 20226 78
rect 20283 42 20290 98
rect 20278 26 20290 42
rect 20215 15 20290 26
rect 20405 98 20480 115
rect 20405 78 20417 98
rect 20405 26 20416 78
rect 20473 42 20480 98
rect 20468 26 20480 42
rect 20405 15 20480 26
rect 20600 98 20675 115
rect 20600 78 20612 98
rect 20600 26 20611 78
rect 20668 42 20675 98
rect 20663 26 20675 42
rect 20600 15 20675 26
rect 20790 98 20865 115
rect 20790 78 20802 98
rect 20790 26 20801 78
rect 20858 42 20865 98
rect 20853 26 20865 42
rect 20790 15 20865 26
rect 20980 98 21055 115
rect 20980 78 20992 98
rect 20980 26 20991 78
rect 21048 42 21055 98
rect 21043 26 21055 42
rect 20980 15 21055 26
rect 21175 98 21250 115
rect 21175 78 21187 98
rect 21175 26 21186 78
rect 21243 42 21250 98
rect 21238 26 21250 42
rect 21175 15 21250 26
rect 21365 98 21440 115
rect 21365 78 21377 98
rect 21365 26 21376 78
rect 21433 42 21440 98
rect 21428 26 21440 42
rect 21365 15 21440 26
rect 21555 98 21630 115
rect 21555 78 21567 98
rect 21555 26 21566 78
rect 21623 42 21630 98
rect 21618 26 21630 42
rect 21555 15 21630 26
rect 21750 98 21825 115
rect 21750 78 21762 98
rect 21750 26 21761 78
rect 21818 42 21825 98
rect 21813 26 21825 42
rect 21750 15 21825 26
rect 8845 -47 11835 -40
rect 8845 -99 9956 -47
rect 10008 -99 10151 -47
rect 10203 -99 10341 -47
rect 10393 -99 10531 -47
rect 10583 -99 10721 -47
rect 10773 -99 10911 -47
rect 10963 -99 11106 -47
rect 11158 -99 11301 -47
rect 11353 -99 11491 -47
rect 11543 -99 11686 -47
rect 11738 -99 11835 -47
rect 8845 -340 11835 -99
rect 12140 -47 12565 -35
rect 12140 -99 12256 -47
rect 12308 -99 12446 -47
rect 12498 -99 12565 -47
rect 8845 -1300 9445 -340
rect 12140 -370 12565 -99
rect 13785 -47 13860 -35
rect 13785 -99 13796 -47
rect 13848 -62 13860 -47
rect 13785 -118 13797 -99
rect 13853 -118 13860 -62
rect 13785 -135 13860 -118
rect 13975 -47 14050 -35
rect 13975 -99 13986 -47
rect 14038 -62 14050 -47
rect 13975 -118 13987 -99
rect 14043 -118 14050 -62
rect 13975 -135 14050 -118
rect 14170 -47 14245 -35
rect 14170 -99 14181 -47
rect 14233 -62 14245 -47
rect 14170 -118 14182 -99
rect 14238 -118 14245 -62
rect 14170 -135 14245 -118
rect 14360 -47 14435 -35
rect 14360 -99 14371 -47
rect 14423 -62 14435 -47
rect 14360 -118 14372 -99
rect 14428 -118 14435 -62
rect 14360 -135 14435 -118
rect 14550 -47 14625 -35
rect 14550 -99 14561 -47
rect 14613 -62 14625 -47
rect 14550 -118 14562 -99
rect 14618 -118 14625 -62
rect 14550 -135 14625 -118
rect 14745 -47 14820 -35
rect 14745 -99 14756 -47
rect 14808 -62 14820 -47
rect 14745 -118 14757 -99
rect 14813 -118 14820 -62
rect 14745 -135 14820 -118
rect 14935 -47 15010 -35
rect 14935 -99 14946 -47
rect 14998 -62 15010 -47
rect 14935 -118 14947 -99
rect 15003 -118 15010 -62
rect 14935 -135 15010 -118
rect 15130 -47 15205 -35
rect 15130 -99 15141 -47
rect 15193 -62 15205 -47
rect 15130 -118 15142 -99
rect 15198 -118 15205 -62
rect 15130 -135 15205 -118
rect 15320 -47 15395 -35
rect 15320 -99 15331 -47
rect 15383 -62 15395 -47
rect 15320 -118 15332 -99
rect 15388 -118 15395 -62
rect 15320 -135 15395 -118
rect 15510 -47 15585 -35
rect 15510 -99 15521 -47
rect 15573 -62 15585 -47
rect 15510 -118 15522 -99
rect 15578 -118 15585 -62
rect 15510 -135 15585 -118
rect 16085 -47 16160 -35
rect 16085 -62 16096 -47
rect 16085 -118 16092 -62
rect 16148 -118 16160 -47
rect 16085 -135 16160 -118
rect 16275 -47 16350 -35
rect 16275 -62 16286 -47
rect 16275 -118 16282 -62
rect 16338 -118 16350 -47
rect 16275 -135 16350 -118
rect 16470 -47 16545 -35
rect 16470 -62 16481 -47
rect 16470 -118 16477 -62
rect 16533 -118 16545 -47
rect 16470 -135 16545 -118
rect 16660 -47 16735 -35
rect 16660 -62 16671 -47
rect 16660 -118 16667 -62
rect 16723 -118 16735 -47
rect 16660 -135 16735 -118
rect 16855 -47 16930 -35
rect 16855 -62 16866 -47
rect 16855 -118 16862 -62
rect 16918 -118 16930 -47
rect 16855 -135 16930 -118
rect 17040 -47 17115 -35
rect 17040 -62 17051 -47
rect 17040 -118 17047 -62
rect 17103 -118 17115 -47
rect 17040 -135 17115 -118
rect 17240 -47 17315 -35
rect 17240 -62 17251 -47
rect 17240 -118 17247 -62
rect 17303 -118 17315 -47
rect 17240 -135 17315 -118
rect 17425 -47 17500 -35
rect 17425 -62 17436 -47
rect 17425 -118 17432 -62
rect 17488 -118 17500 -47
rect 17425 -135 17500 -118
rect 17620 -47 17695 -35
rect 17620 -62 17631 -47
rect 17620 -118 17627 -62
rect 17683 -118 17695 -47
rect 17620 -135 17695 -118
rect 17815 -47 17890 -35
rect 17815 -62 17826 -47
rect 17815 -118 17822 -62
rect 17878 -118 17890 -47
rect 17815 -135 17890 -118
rect 18000 -47 18075 -35
rect 18000 -62 18011 -47
rect 18000 -118 18007 -62
rect 18063 -118 18075 -47
rect 18000 -135 18075 -118
rect 18195 -47 18270 -35
rect 18195 -62 18206 -47
rect 18195 -118 18202 -62
rect 18258 -118 18270 -47
rect 18195 -135 18270 -118
rect 18385 -47 18460 -35
rect 18385 -62 18396 -47
rect 18385 -118 18392 -62
rect 18448 -118 18460 -47
rect 18385 -135 18460 -118
rect 18580 -47 18655 -35
rect 18580 -62 18591 -47
rect 18580 -118 18587 -62
rect 18643 -118 18655 -47
rect 18580 -135 18655 -118
rect 18770 -47 18845 -35
rect 18770 -62 18781 -47
rect 18770 -118 18777 -62
rect 18833 -118 18845 -47
rect 18770 -135 18845 -118
rect 18965 -47 19040 -35
rect 18965 -62 18976 -47
rect 18965 -118 18972 -62
rect 19028 -118 19040 -47
rect 18965 -135 19040 -118
rect 19155 -47 19230 -35
rect 19155 -62 19166 -47
rect 19155 -118 19162 -62
rect 19218 -118 19230 -47
rect 19155 -135 19230 -118
rect 19350 -47 19425 -35
rect 19350 -62 19361 -47
rect 19350 -118 19357 -62
rect 19413 -118 19425 -47
rect 19350 -135 19425 -118
rect 19540 -47 19615 -35
rect 19540 -62 19551 -47
rect 19540 -118 19547 -62
rect 19603 -118 19615 -47
rect 19540 -135 19615 -118
rect 19735 -47 19810 -35
rect 19735 -62 19746 -47
rect 19735 -118 19742 -62
rect 19798 -118 19810 -47
rect 19735 -135 19810 -118
rect 19925 -47 20000 -35
rect 19925 -62 19936 -47
rect 19925 -118 19932 -62
rect 19988 -118 20000 -47
rect 19925 -135 20000 -118
rect 20115 -47 20190 -35
rect 20115 -62 20126 -47
rect 20115 -118 20122 -62
rect 20178 -118 20190 -47
rect 20115 -135 20190 -118
rect 20310 -47 20385 -35
rect 20310 -62 20321 -47
rect 20310 -118 20317 -62
rect 20373 -118 20385 -47
rect 20310 -135 20385 -118
rect 20500 -47 20575 -35
rect 20500 -62 20511 -47
rect 20500 -118 20507 -62
rect 20563 -118 20575 -47
rect 20500 -135 20575 -118
rect 20695 -47 20770 -35
rect 20695 -62 20706 -47
rect 20695 -118 20702 -62
rect 20758 -118 20770 -47
rect 20695 -135 20770 -118
rect 20885 -47 20960 -35
rect 20885 -62 20896 -47
rect 20885 -118 20892 -62
rect 20948 -118 20960 -47
rect 20885 -135 20960 -118
rect 21075 -47 21150 -35
rect 21075 -62 21086 -47
rect 21075 -118 21082 -62
rect 21138 -118 21150 -47
rect 21075 -135 21150 -118
rect 21270 -47 21345 -35
rect 21270 -62 21281 -47
rect 21270 -118 21277 -62
rect 21333 -118 21345 -47
rect 21270 -135 21345 -118
rect 21460 -47 21535 -35
rect 21460 -62 21471 -47
rect 21460 -118 21467 -62
rect 21523 -118 21535 -47
rect 21460 -135 21535 -118
rect 21650 -47 21725 -35
rect 21650 -62 21661 -47
rect 21650 -118 21657 -62
rect 21713 -118 21725 -47
rect 21650 -135 21725 -118
rect 13515 -157 13590 -145
rect 13515 -209 13526 -157
rect 13578 -209 13590 -157
rect 13515 -370 13590 -209
rect 12140 -440 13590 -370
rect 10190 -565 10615 -520
rect 10190 -587 10216 -565
rect 10588 -587 10615 -565
rect 10190 -1043 10214 -587
rect 10590 -1043 10615 -587
rect 10190 -1065 10216 -1043
rect 10588 -1065 10615 -1043
rect 10190 -1090 10615 -1065
rect 12140 -558 12565 -440
rect 12140 -1058 12169 -558
rect 12541 -1058 12565 -558
rect 12140 -1090 12565 -1058
rect 13725 -570 14165 -520
rect 13725 -600 13756 -570
rect 14128 -600 14165 -570
rect 13725 -1616 13754 -600
rect 14130 -1616 14165 -600
rect 13725 -1646 13756 -1616
rect 14128 -1646 14165 -1616
rect 13725 -1675 14165 -1646
rect 17435 -572 17870 -530
rect 17435 -602 17466 -572
rect 17838 -602 17870 -572
rect 17435 -1618 17464 -602
rect 17840 -1618 17870 -602
rect 17435 -1648 17466 -1618
rect 17838 -1648 17870 -1618
rect 17435 -1675 17870 -1648
<< via2 >>
rect 10219 1227 10221 1683
rect 10221 1227 10593 1683
rect 10593 1227 10595 1683
rect 13742 1227 13744 2243
rect 13744 1227 14116 2243
rect 14116 1227 14118 2243
rect 17459 1227 17461 2243
rect 17461 1227 17833 2243
rect 17833 1227 17835 2243
rect 13797 738 13853 758
rect 13797 702 13848 738
rect 13848 702 13853 738
rect 13987 738 14043 758
rect 13987 702 14038 738
rect 14038 702 14043 738
rect 14182 738 14238 758
rect 14182 702 14233 738
rect 14233 702 14238 738
rect 14372 738 14428 758
rect 14372 702 14423 738
rect 14423 702 14428 738
rect 14562 738 14618 758
rect 14562 702 14613 738
rect 14613 702 14618 738
rect 14757 738 14813 758
rect 14757 702 14808 738
rect 14808 702 14813 738
rect 14947 738 15003 758
rect 14947 702 14998 738
rect 14998 702 15003 738
rect 15142 738 15198 758
rect 15142 702 15193 738
rect 15193 702 15198 738
rect 15332 738 15388 758
rect 15332 702 15383 738
rect 15383 702 15388 738
rect 15522 738 15578 758
rect 15522 702 15573 738
rect 15573 702 15578 738
rect 16092 738 16148 758
rect 16092 702 16096 738
rect 16096 702 16148 738
rect 16282 738 16338 758
rect 16282 702 16286 738
rect 16286 702 16338 738
rect 16477 738 16533 758
rect 16477 702 16481 738
rect 16481 702 16533 738
rect 16667 738 16723 758
rect 16667 702 16671 738
rect 16671 702 16723 738
rect 16862 738 16918 758
rect 16862 702 16866 738
rect 16866 702 16918 738
rect 17047 738 17103 758
rect 17047 702 17051 738
rect 17051 702 17103 738
rect 17247 738 17303 758
rect 17247 702 17251 738
rect 17251 702 17303 738
rect 17432 738 17488 758
rect 17432 702 17436 738
rect 17436 702 17488 738
rect 17627 738 17683 758
rect 17627 702 17631 738
rect 17631 702 17683 738
rect 17822 738 17878 758
rect 17822 702 17826 738
rect 17826 702 17878 738
rect 18007 738 18063 758
rect 18007 702 18011 738
rect 18011 702 18063 738
rect 18202 738 18258 758
rect 18202 702 18206 738
rect 18206 702 18258 738
rect 18392 738 18448 758
rect 18392 702 18396 738
rect 18396 702 18448 738
rect 18587 738 18643 758
rect 18587 702 18591 738
rect 18591 702 18643 738
rect 18777 738 18833 758
rect 18777 702 18781 738
rect 18781 702 18833 738
rect 18972 738 19028 758
rect 18972 702 18976 738
rect 18976 702 19028 738
rect 19162 738 19218 758
rect 19162 702 19166 738
rect 19166 702 19218 738
rect 19357 738 19413 758
rect 19357 702 19361 738
rect 19361 702 19413 738
rect 19547 738 19603 758
rect 19547 702 19551 738
rect 19551 702 19603 738
rect 19742 738 19798 758
rect 19742 702 19746 738
rect 19746 702 19798 738
rect 19932 738 19988 758
rect 19932 702 19936 738
rect 19936 702 19988 738
rect 20122 738 20178 758
rect 20122 702 20126 738
rect 20126 702 20178 738
rect 20317 738 20373 758
rect 20317 702 20321 738
rect 20321 702 20373 738
rect 20507 738 20563 758
rect 20507 702 20511 738
rect 20511 702 20563 738
rect 20702 738 20758 758
rect 20702 702 20706 738
rect 20706 702 20758 738
rect 20892 738 20948 758
rect 20892 702 20896 738
rect 20896 702 20948 738
rect 21082 738 21138 758
rect 21082 702 21086 738
rect 21086 702 21138 738
rect 21277 738 21333 758
rect 21277 702 21281 738
rect 21281 702 21333 738
rect 21467 738 21523 758
rect 21467 702 21471 738
rect 21471 702 21523 738
rect 21657 738 21713 758
rect 21657 702 21661 738
rect 21661 702 21713 738
rect 13702 561 13753 598
rect 13753 561 13758 598
rect 13702 542 13758 561
rect 13892 561 13943 598
rect 13943 561 13948 598
rect 13892 542 13948 561
rect 14087 561 14138 598
rect 14138 561 14143 598
rect 14087 542 14143 561
rect 14277 561 14328 598
rect 14328 561 14333 598
rect 14277 542 14333 561
rect 14472 561 14523 598
rect 14523 561 14528 598
rect 14472 542 14528 561
rect 14657 561 14708 598
rect 14708 561 14713 598
rect 14657 542 14713 561
rect 14852 561 14903 598
rect 14903 561 14908 598
rect 14852 542 14908 561
rect 15042 561 15093 598
rect 15093 561 15098 598
rect 15042 542 15098 561
rect 15237 561 15288 598
rect 15288 561 15293 598
rect 15237 542 15293 561
rect 15427 561 15478 598
rect 15478 561 15483 598
rect 15427 542 15483 561
rect 15622 561 15673 598
rect 15673 561 15678 598
rect 15622 542 15678 561
rect 15997 561 16048 598
rect 16048 561 16053 598
rect 15997 542 16053 561
rect 16187 561 16238 598
rect 16238 561 16243 598
rect 16187 542 16243 561
rect 16382 561 16433 598
rect 16433 561 16438 598
rect 16382 542 16438 561
rect 16577 561 16628 598
rect 16628 561 16633 598
rect 16577 542 16633 561
rect 16767 561 16818 598
rect 16818 561 16823 598
rect 16767 542 16823 561
rect 16962 561 17013 598
rect 17013 561 17018 598
rect 16962 542 17018 561
rect 17152 561 17203 598
rect 17203 561 17208 598
rect 17152 542 17208 561
rect 17347 561 17398 598
rect 17398 561 17403 598
rect 17347 542 17403 561
rect 17537 561 17588 598
rect 17588 561 17593 598
rect 17537 542 17593 561
rect 17727 561 17778 598
rect 17778 561 17783 598
rect 17727 542 17783 561
rect 17922 561 17973 598
rect 17973 561 17978 598
rect 17922 542 17978 561
rect 18112 561 18163 598
rect 18163 561 18168 598
rect 18112 542 18168 561
rect 18307 561 18358 598
rect 18358 561 18363 598
rect 18307 542 18363 561
rect 18497 561 18548 598
rect 18548 561 18553 598
rect 18497 542 18553 561
rect 18687 561 18738 598
rect 18738 561 18743 598
rect 18687 542 18743 561
rect 18882 561 18933 598
rect 18933 561 18938 598
rect 18882 542 18938 561
rect 19072 561 19123 598
rect 19123 561 19128 598
rect 19072 542 19128 561
rect 19267 561 19318 598
rect 19318 561 19323 598
rect 19267 542 19323 561
rect 19457 561 19508 598
rect 19508 561 19513 598
rect 19457 542 19513 561
rect 19647 561 19698 598
rect 19698 561 19703 598
rect 19647 542 19703 561
rect 19842 561 19893 598
rect 19893 561 19898 598
rect 19842 542 19898 561
rect 20032 561 20083 598
rect 20083 561 20088 598
rect 20032 542 20088 561
rect 20227 561 20278 598
rect 20278 561 20283 598
rect 20227 542 20283 561
rect 20417 561 20468 598
rect 20468 561 20473 598
rect 20417 542 20473 561
rect 20612 561 20663 598
rect 20663 561 20668 598
rect 20612 542 20668 561
rect 20802 561 20853 598
rect 20853 561 20858 598
rect 20802 542 20858 561
rect 20992 561 21043 598
rect 21043 561 21048 598
rect 20992 542 21048 561
rect 21187 561 21238 598
rect 21238 561 21243 598
rect 21187 542 21243 561
rect 21377 561 21428 598
rect 21428 561 21433 598
rect 21377 542 21433 561
rect 21567 561 21618 598
rect 21618 561 21623 598
rect 21567 542 21623 561
rect 21762 561 21813 598
rect 21813 561 21818 598
rect 21762 542 21818 561
rect 13702 78 13758 98
rect 13702 42 13753 78
rect 13753 42 13758 78
rect 13892 78 13948 98
rect 13892 42 13943 78
rect 13943 42 13948 78
rect 14087 78 14143 98
rect 14087 42 14138 78
rect 14138 42 14143 78
rect 14277 78 14333 98
rect 14277 42 14328 78
rect 14328 42 14333 78
rect 14472 78 14528 98
rect 14472 42 14523 78
rect 14523 42 14528 78
rect 14657 78 14713 98
rect 14657 42 14708 78
rect 14708 42 14713 78
rect 14852 78 14908 98
rect 14852 42 14903 78
rect 14903 42 14908 78
rect 15042 78 15098 98
rect 15042 42 15093 78
rect 15093 42 15098 78
rect 15237 78 15293 98
rect 15237 42 15288 78
rect 15288 42 15293 78
rect 15427 78 15483 98
rect 15427 42 15478 78
rect 15478 42 15483 78
rect 15622 78 15678 98
rect 15622 42 15673 78
rect 15673 42 15678 78
rect 15997 78 16053 98
rect 15997 42 16048 78
rect 16048 42 16053 78
rect 16187 78 16243 98
rect 16187 42 16238 78
rect 16238 42 16243 78
rect 16382 78 16438 98
rect 16382 42 16433 78
rect 16433 42 16438 78
rect 16577 78 16633 98
rect 16577 42 16628 78
rect 16628 42 16633 78
rect 16767 78 16823 98
rect 16767 42 16818 78
rect 16818 42 16823 78
rect 16962 78 17018 98
rect 16962 42 17013 78
rect 17013 42 17018 78
rect 17152 78 17208 98
rect 17152 42 17203 78
rect 17203 42 17208 78
rect 17347 78 17403 98
rect 17347 42 17398 78
rect 17398 42 17403 78
rect 17537 78 17593 98
rect 17537 42 17588 78
rect 17588 42 17593 78
rect 17727 78 17783 98
rect 17727 42 17778 78
rect 17778 42 17783 78
rect 17922 78 17978 98
rect 17922 42 17973 78
rect 17973 42 17978 78
rect 18112 78 18168 98
rect 18112 42 18163 78
rect 18163 42 18168 78
rect 18307 78 18363 98
rect 18307 42 18358 78
rect 18358 42 18363 78
rect 18497 78 18553 98
rect 18497 42 18548 78
rect 18548 42 18553 78
rect 18687 78 18743 98
rect 18687 42 18738 78
rect 18738 42 18743 78
rect 18882 78 18938 98
rect 18882 42 18933 78
rect 18933 42 18938 78
rect 19072 78 19128 98
rect 19072 42 19123 78
rect 19123 42 19128 78
rect 19267 78 19323 98
rect 19267 42 19318 78
rect 19318 42 19323 78
rect 19457 78 19513 98
rect 19457 42 19508 78
rect 19508 42 19513 78
rect 19647 78 19703 98
rect 19647 42 19698 78
rect 19698 42 19703 78
rect 19842 78 19898 98
rect 19842 42 19893 78
rect 19893 42 19898 78
rect 20032 78 20088 98
rect 20032 42 20083 78
rect 20083 42 20088 78
rect 20227 78 20283 98
rect 20227 42 20278 78
rect 20278 42 20283 78
rect 20417 78 20473 98
rect 20417 42 20468 78
rect 20468 42 20473 78
rect 20612 78 20668 98
rect 20612 42 20663 78
rect 20663 42 20668 78
rect 20802 78 20858 98
rect 20802 42 20853 78
rect 20853 42 20858 78
rect 20992 78 21048 98
rect 20992 42 21043 78
rect 21043 42 21048 78
rect 21187 78 21243 98
rect 21187 42 21238 78
rect 21238 42 21243 78
rect 21377 78 21433 98
rect 21377 42 21428 78
rect 21428 42 21433 78
rect 21567 78 21623 98
rect 21567 42 21618 78
rect 21618 42 21623 78
rect 21762 78 21818 98
rect 21762 42 21813 78
rect 21813 42 21818 78
rect 13797 -99 13848 -62
rect 13848 -99 13853 -62
rect 13797 -118 13853 -99
rect 13987 -99 14038 -62
rect 14038 -99 14043 -62
rect 13987 -118 14043 -99
rect 14182 -99 14233 -62
rect 14233 -99 14238 -62
rect 14182 -118 14238 -99
rect 14372 -99 14423 -62
rect 14423 -99 14428 -62
rect 14372 -118 14428 -99
rect 14562 -99 14613 -62
rect 14613 -99 14618 -62
rect 14562 -118 14618 -99
rect 14757 -99 14808 -62
rect 14808 -99 14813 -62
rect 14757 -118 14813 -99
rect 14947 -99 14998 -62
rect 14998 -99 15003 -62
rect 14947 -118 15003 -99
rect 15142 -99 15193 -62
rect 15193 -99 15198 -62
rect 15142 -118 15198 -99
rect 15332 -99 15383 -62
rect 15383 -99 15388 -62
rect 15332 -118 15388 -99
rect 15522 -99 15573 -62
rect 15573 -99 15578 -62
rect 15522 -118 15578 -99
rect 16092 -99 16096 -62
rect 16096 -99 16148 -62
rect 16092 -118 16148 -99
rect 16282 -99 16286 -62
rect 16286 -99 16338 -62
rect 16282 -118 16338 -99
rect 16477 -99 16481 -62
rect 16481 -99 16533 -62
rect 16477 -118 16533 -99
rect 16667 -99 16671 -62
rect 16671 -99 16723 -62
rect 16667 -118 16723 -99
rect 16862 -99 16866 -62
rect 16866 -99 16918 -62
rect 16862 -118 16918 -99
rect 17047 -99 17051 -62
rect 17051 -99 17103 -62
rect 17047 -118 17103 -99
rect 17247 -99 17251 -62
rect 17251 -99 17303 -62
rect 17247 -118 17303 -99
rect 17432 -99 17436 -62
rect 17436 -99 17488 -62
rect 17432 -118 17488 -99
rect 17627 -99 17631 -62
rect 17631 -99 17683 -62
rect 17627 -118 17683 -99
rect 17822 -99 17826 -62
rect 17826 -99 17878 -62
rect 17822 -118 17878 -99
rect 18007 -99 18011 -62
rect 18011 -99 18063 -62
rect 18007 -118 18063 -99
rect 18202 -99 18206 -62
rect 18206 -99 18258 -62
rect 18202 -118 18258 -99
rect 18392 -99 18396 -62
rect 18396 -99 18448 -62
rect 18392 -118 18448 -99
rect 18587 -99 18591 -62
rect 18591 -99 18643 -62
rect 18587 -118 18643 -99
rect 18777 -99 18781 -62
rect 18781 -99 18833 -62
rect 18777 -118 18833 -99
rect 18972 -99 18976 -62
rect 18976 -99 19028 -62
rect 18972 -118 19028 -99
rect 19162 -99 19166 -62
rect 19166 -99 19218 -62
rect 19162 -118 19218 -99
rect 19357 -99 19361 -62
rect 19361 -99 19413 -62
rect 19357 -118 19413 -99
rect 19547 -99 19551 -62
rect 19551 -99 19603 -62
rect 19547 -118 19603 -99
rect 19742 -99 19746 -62
rect 19746 -99 19798 -62
rect 19742 -118 19798 -99
rect 19932 -99 19936 -62
rect 19936 -99 19988 -62
rect 19932 -118 19988 -99
rect 20122 -99 20126 -62
rect 20126 -99 20178 -62
rect 20122 -118 20178 -99
rect 20317 -99 20321 -62
rect 20321 -99 20373 -62
rect 20317 -118 20373 -99
rect 20507 -99 20511 -62
rect 20511 -99 20563 -62
rect 20507 -118 20563 -99
rect 20702 -99 20706 -62
rect 20706 -99 20758 -62
rect 20702 -118 20758 -99
rect 20892 -99 20896 -62
rect 20896 -99 20948 -62
rect 20892 -118 20948 -99
rect 21082 -99 21086 -62
rect 21086 -99 21138 -62
rect 21082 -118 21138 -99
rect 21277 -99 21281 -62
rect 21281 -99 21333 -62
rect 21277 -118 21333 -99
rect 21467 -99 21471 -62
rect 21471 -99 21523 -62
rect 21467 -118 21523 -99
rect 21657 -99 21661 -62
rect 21661 -99 21713 -62
rect 21657 -118 21713 -99
rect 10214 -1043 10216 -587
rect 10216 -1043 10588 -587
rect 10588 -1043 10590 -587
rect 13754 -1616 13756 -600
rect 13756 -1616 14128 -600
rect 14128 -1616 14130 -600
rect 17464 -1618 17466 -602
rect 17466 -1618 17838 -602
rect 17838 -1618 17840 -602
<< metal3 >>
rect 13725 2320 14160 2475
rect 13715 2243 14160 2320
rect 10190 1683 10640 1735
rect 10190 1227 10219 1683
rect 10595 1227 10640 1683
rect 10190 -587 10640 1227
rect 13715 1227 13742 2243
rect 14118 2040 14160 2243
rect 17435 2247 17870 2310
rect 14118 1227 14150 2040
rect 13715 1090 14150 1227
rect 17435 1223 17455 2247
rect 17839 1223 17870 2247
rect 17435 1165 17870 1223
rect 13715 758 15710 1090
rect 13715 745 13797 758
rect 13785 702 13797 745
rect 13853 702 13987 758
rect 14043 702 14182 758
rect 14238 702 14372 758
rect 14428 702 14562 758
rect 14618 702 14757 758
rect 14813 702 14947 758
rect 15003 702 15142 758
rect 15198 702 15332 758
rect 15388 702 15522 758
rect 15578 702 15710 758
rect 13785 685 15710 702
rect 15980 765 22825 1100
rect 15980 758 21820 765
rect 15980 702 16092 758
rect 16148 702 16282 758
rect 16338 702 16477 758
rect 16533 702 16667 758
rect 16723 702 16862 758
rect 16918 702 17047 758
rect 17103 702 17247 758
rect 17303 702 17432 758
rect 17488 702 17627 758
rect 17683 702 17822 758
rect 17878 702 18007 758
rect 18063 702 18202 758
rect 18258 702 18392 758
rect 18448 702 18587 758
rect 18643 702 18777 758
rect 18833 702 18972 758
rect 19028 702 19162 758
rect 19218 702 19357 758
rect 19413 702 19547 758
rect 19603 702 19742 758
rect 19798 702 19932 758
rect 19988 702 20122 758
rect 20178 702 20317 758
rect 20373 702 20507 758
rect 20563 702 20702 758
rect 20758 702 20892 758
rect 20948 702 21082 758
rect 21138 702 21277 758
rect 21333 702 21467 758
rect 21523 702 21657 758
rect 21713 702 21820 758
rect 15980 685 21820 702
rect 13680 598 21825 615
rect 13680 542 13702 598
rect 13758 542 13892 598
rect 13948 542 14087 598
rect 14143 542 14277 598
rect 14333 542 14472 598
rect 14528 542 14657 598
rect 14713 542 14852 598
rect 14908 542 15042 598
rect 15098 542 15237 598
rect 15293 542 15427 598
rect 15483 542 15622 598
rect 15678 542 15997 598
rect 16053 542 16187 598
rect 16243 542 16382 598
rect 16438 542 16577 598
rect 16633 542 16767 598
rect 16823 542 16962 598
rect 17018 542 17152 598
rect 17208 542 17347 598
rect 17403 542 17537 598
rect 17593 542 17727 598
rect 17783 542 17922 598
rect 17978 542 18112 598
rect 18168 542 18307 598
rect 18363 542 18497 598
rect 18553 542 18687 598
rect 18743 542 18882 598
rect 18938 542 19072 598
rect 19128 542 19267 598
rect 19323 542 19457 598
rect 19513 542 19647 598
rect 19703 542 19842 598
rect 19898 542 20032 598
rect 20088 542 20227 598
rect 20283 542 20417 598
rect 20473 542 20612 598
rect 20668 542 20802 598
rect 20858 542 20992 598
rect 21048 542 21187 598
rect 21243 542 21377 598
rect 21433 542 21567 598
rect 21623 542 21762 598
rect 21818 542 21825 598
rect 13680 98 21825 542
rect 13680 42 13702 98
rect 13758 42 13892 98
rect 13948 42 14087 98
rect 14143 42 14277 98
rect 14333 42 14472 98
rect 14528 42 14657 98
rect 14713 42 14852 98
rect 14908 42 15042 98
rect 15098 42 15237 98
rect 15293 42 15427 98
rect 15483 42 15622 98
rect 15678 42 15997 98
rect 16053 42 16187 98
rect 16243 42 16382 98
rect 16438 42 16577 98
rect 16633 42 16767 98
rect 16823 42 16962 98
rect 17018 42 17152 98
rect 17208 42 17347 98
rect 17403 42 17537 98
rect 17593 42 17727 98
rect 17783 42 17922 98
rect 17978 42 18112 98
rect 18168 42 18307 98
rect 18363 42 18497 98
rect 18553 42 18687 98
rect 18743 42 18882 98
rect 18938 42 19072 98
rect 19128 42 19267 98
rect 19323 42 19457 98
rect 19513 42 19647 98
rect 19703 42 19842 98
rect 19898 42 20032 98
rect 20088 42 20227 98
rect 20283 42 20417 98
rect 20473 42 20612 98
rect 20668 42 20802 98
rect 20858 42 20992 98
rect 21048 42 21187 98
rect 21243 42 21377 98
rect 21433 42 21567 98
rect 21623 42 21762 98
rect 21818 42 21825 98
rect 13680 25 21825 42
rect 22025 -45 22825 765
rect 10190 -1043 10214 -587
rect 10590 -1043 10640 -587
rect 10190 -1275 10640 -1043
rect 13725 -62 15710 -45
rect 13725 -118 13797 -62
rect 13853 -118 13987 -62
rect 14043 -118 14182 -62
rect 14238 -118 14372 -62
rect 14428 -118 14562 -62
rect 14618 -118 14757 -62
rect 14813 -118 14947 -62
rect 15003 -118 15142 -62
rect 15198 -118 15332 -62
rect 15388 -118 15522 -62
rect 15578 -118 15710 -62
rect 13725 -455 15710 -118
rect 15980 -62 22825 -45
rect 15980 -118 16092 -62
rect 16148 -118 16282 -62
rect 16338 -118 16477 -62
rect 16533 -118 16667 -62
rect 16723 -118 16862 -62
rect 16918 -118 17047 -62
rect 17103 -118 17247 -62
rect 17303 -118 17432 -62
rect 17488 -118 17627 -62
rect 17683 -118 17822 -62
rect 17878 -118 18007 -62
rect 18063 -118 18202 -62
rect 18258 -118 18392 -62
rect 18448 -118 18587 -62
rect 18643 -118 18777 -62
rect 18833 -118 18972 -62
rect 19028 -118 19162 -62
rect 19218 -118 19357 -62
rect 19413 -118 19547 -62
rect 19603 -118 19742 -62
rect 19798 -118 19932 -62
rect 19988 -118 20122 -62
rect 20178 -118 20317 -62
rect 20373 -118 20507 -62
rect 20563 -118 20702 -62
rect 20758 -118 20892 -62
rect 20948 -118 21082 -62
rect 21138 -118 21277 -62
rect 21333 -118 21467 -62
rect 21523 -118 21657 -62
rect 21713 -118 22825 -62
rect 15980 -455 22825 -118
rect 13725 -600 14160 -455
rect 13725 -1616 13754 -600
rect 14130 -1430 14160 -600
rect 17435 -598 17870 -530
rect 14130 -1616 14165 -1430
rect 13725 -1680 14165 -1616
rect 17435 -1622 17460 -598
rect 17844 -1622 17870 -598
rect 17435 -1675 17870 -1622
rect 13730 -1865 14165 -1680
rect 22025 -1795 22825 -455
<< via3 >>
rect 17455 2243 17839 2247
rect 17455 1227 17459 2243
rect 17459 1227 17835 2243
rect 17835 1227 17839 2243
rect 17455 1223 17839 1227
rect 17460 -602 17844 -598
rect 17460 -1618 17464 -602
rect 17464 -1618 17840 -602
rect 17840 -1618 17844 -602
rect 17460 -1622 17844 -1618
<< metal4 >>
rect 17435 2247 18025 2310
rect 17435 1223 17455 2247
rect 17839 1223 18025 2247
rect 17435 -598 18025 1223
rect 17435 -1622 17460 -598
rect 17844 -1622 18025 -598
rect 17435 -1675 18025 -1622
rect 17440 -1680 18025 -1675
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM1
timestamp 1663011646
transform 1 0 10847 0 -1 650
box -1117 -300 1117 300
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM2
timestamp 1663011646
transform 1 0 10847 0 1 -10
box -1117 -300 1117 300
use sky130_fd_pr__nfet_01v8_lvt_LELFGX  XM3
timestamp 1663011646
transform 1 0 18902 0 1 650
box -3037 -300 3037 300
use sky130_fd_pr__nfet_01v8_lvt_LELFGX  XM4
timestamp 1663011646
transform 1 0 18902 0 1 -10
box -3037 -300 3037 300
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM32
timestamp 1663011646
transform 1 0 14687 0 1 650
box -1117 -300 1117 300
use sky130_fd_pr__nfet_01v8_lvt_YTLFGX  XM33
timestamp 1663011646
transform 1 0 14687 0 -1 -10
box -1117 -300 1117 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM42
timestamp 1663011646
transform 1 0 12379 0 -1 650
box -349 -300 349 300
use sky130_fd_pr__nfet_01v8_lvt_HNLS5R  XM43
timestamp 1663011646
transform 1 0 12379 0 1 -10
box -349 -300 349 300
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR1
timestamp 1663011646
transform 0 1 11383 -1 0 1451
box -441 -1348 441 1348
use sky130_fd_pr__res_high_po_2p85_P79JE3  XR2
timestamp 1663011646
transform 0 1 11380 -1 0 -807
box -441 -1348 441 1348
use sky130_fd_pr__res_high_po_5p73_W59YBA  XR3
timestamp 1663011646
transform 0 1 15798 -1 0 -1101
box -729 -2228 729 2228
use sky130_fd_pr__res_high_po_5p73_W59YBA  XR29
timestamp 1663011646
transform 0 1 15798 -1 0 1739
box -729 -2228 729 2228
<< labels >>
rlabel metal1 s 11925 -1260 11975 830 4 BIAS
port 1 nsew
rlabel metal2 s 8845 -1300 9445 980 4 GND
port 2 nsew
rlabel metal3 s 10190 -1275 10640 -1080 4 VDD
port 3 nsew
rlabel metal1 s 12900 -1255 12955 175 4 INB
port 4 nsew
rlabel metal1 s 13365 -1260 13415 520 4 INA
port 5 nsew
rlabel metal3 s 22025 -1795 22825 -240 4 GND
port 2 nsew
rlabel metal4 s 17440 -1680 18025 2310 4 VDD
port 3 nsew
rlabel metal1 s 15855 -1840 15905 830 4 BIAS
port 1 nsew
rlabel locali s 12675 1830 13610 1870 4 SUB
port 6 nsew
rlabel metal3 s 13725 2280 14160 2475 4 OUTA
port 7 nsew
rlabel metal3 s 13730 -1865 14165 -1655 4 OUTB
port 8 nsew
<< end >>
