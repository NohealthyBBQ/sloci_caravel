magic
tech sky130A
magscale 1 2
timestamp 1666262589
<< metal1 >>
rect 491912 626638 491922 626694
rect 491978 626638 491988 626694
rect 491911 626492 491921 626548
rect 491977 626492 491987 626548
rect 515895 569455 515905 569669
rect 516059 569455 516069 569669
rect 491495 565936 491505 566596
rect 491689 565936 491699 566596
rect 513768 559273 513778 559279
rect 513447 559222 513778 559273
rect 513768 559215 513778 559222
rect 513842 559215 513852 559279
rect 496803 559068 496813 559132
rect 496877 559068 496887 559132
rect 444689 450571 444699 450765
rect 444321 450566 444699 450571
rect 445166 450566 445176 450765
rect 444321 449797 445060 450566
rect 444321 418953 445054 449797
rect 443471 412049 443481 412101
rect 443533 412049 443543 412101
rect 443471 411908 443481 411960
rect 443533 411908 443543 411960
rect 467461 355277 467471 355425
rect 467538 355277 467548 355425
rect 443140 352045 443150 352473
rect 443254 352045 443264 352473
rect 473198 345598 473292 345618
rect 473198 345534 473216 345598
rect 473280 345534 473292 345598
rect 473198 344683 473292 345534
rect 465142 344634 473292 344683
rect 465142 344633 473258 344634
rect 448364 344480 448374 344544
rect 448438 344480 448448 344544
<< via1 >>
rect 491922 626638 491978 626694
rect 491921 626492 491977 626548
rect 515905 569455 516059 569669
rect 491505 565936 491689 566596
rect 513778 559215 513842 559279
rect 496813 559068 496877 559132
rect 444699 450566 445166 450765
rect 443481 412049 443533 412101
rect 443481 411908 443533 411960
rect 467471 355277 467538 355425
rect 443150 352045 443254 352473
rect 473216 345534 473280 345598
rect 448374 344480 448438 344544
<< metal2 >>
rect 493920 633980 494520 633990
rect 493920 633350 494520 633360
rect 494067 632872 494235 633350
rect 491640 626706 491767 626707
rect 491640 626694 491995 626706
rect 491640 626689 491922 626694
rect 491640 626633 491662 626689
rect 491718 626638 491922 626689
rect 491978 626638 491995 626694
rect 491718 626633 491995 626638
rect 491640 626622 491995 626633
rect 491644 626548 491992 626560
rect 491644 626545 491921 626548
rect 491644 626489 491656 626545
rect 491712 626492 491921 626545
rect 491977 626492 491992 626548
rect 491712 626489 491992 626492
rect 491644 626476 491992 626489
rect 491644 626475 491771 626476
rect 486048 595121 487425 595433
rect 486048 594419 486464 595121
rect 487165 594419 487425 595121
rect 486048 559030 487425 594419
rect 515905 569669 516059 569679
rect 515905 569445 516059 569455
rect 491505 566596 491689 566606
rect 491505 565926 491689 565936
rect 513760 559279 513877 559292
rect 513760 559215 513778 559279
rect 513842 559215 513877 559279
rect 513760 559204 513877 559215
rect 496792 559132 496908 559142
rect 496792 559068 496813 559132
rect 496877 559068 496908 559132
rect 496792 559054 496908 559068
rect 486048 557812 486191 559030
rect 487334 557812 487425 559030
rect 486048 557650 487425 557812
rect 446144 453586 461576 453594
rect 446098 453584 461576 453586
rect 446098 453574 446144 453584
rect 445625 451623 446144 453574
rect 445625 451613 461576 451623
rect 444699 450765 445166 450775
rect 444699 450556 445166 450566
rect 445625 418319 446282 451613
rect 403648 412519 403740 412529
rect 403740 412425 443633 412476
rect 403648 412424 443633 412425
rect 403648 412415 403740 412424
rect 443481 412101 443535 412424
rect 443533 412093 443535 412101
rect 443481 412039 443533 412049
rect 403659 411980 403751 411990
rect 403505 411908 403659 411960
rect 443481 411960 443533 411970
rect 403751 411908 443481 411960
rect 443481 411898 443533 411908
rect 403659 411876 403751 411886
rect 467471 355425 467538 355435
rect 467471 355267 467538 355277
rect 443150 352473 443254 352483
rect 443150 352035 443254 352045
rect 473196 345598 473384 345624
rect 473196 345534 473216 345598
rect 473280 345534 473384 345598
rect 473196 345519 473384 345534
rect 448355 344544 448491 344559
rect 448355 344480 448374 344544
rect 448438 344480 448491 344544
rect 448355 344464 448491 344480
<< via2 >>
rect 493920 633360 494520 633980
rect 491662 626633 491718 626689
rect 491656 626489 491712 626545
rect 486464 594419 487165 595121
rect 515905 569455 516059 569669
rect 491505 565936 491689 566596
rect 513778 559215 513842 559279
rect 496813 559068 496877 559132
rect 486191 557812 487334 559030
rect 446144 451623 461576 453584
rect 444699 450566 445166 450765
rect 403648 412425 403740 412519
rect 403659 411886 403751 411980
rect 467471 355277 467538 355425
rect 443150 352045 443254 352473
rect 473216 345534 473280 345598
rect 448374 344480 448438 344544
<< metal3 >>
rect 465334 702380 470924 706352
rect 465334 701598 474059 702380
rect 465370 700807 474059 701598
rect 477386 700807 477803 702380
rect 510002 702246 525998 702538
rect 566570 702380 571314 702382
rect 536597 702282 571314 702380
rect 465370 700584 477803 700807
rect 510000 702000 526000 702246
rect 510000 694000 511000 702000
rect 525000 694000 526000 702000
rect 536597 702106 571317 702282
rect 536597 699875 537573 702106
rect 540501 699875 571317 702106
rect 536597 699317 571317 699875
rect 510000 693000 526000 694000
rect 582224 682863 582500 682892
rect 547752 681190 582500 682863
rect 547752 678122 548589 681190
rect 551656 678122 582500 681190
rect 547752 677972 582500 678122
rect 547752 677425 582490 677972
rect 582248 644600 582858 644604
rect 570200 643000 582858 644600
rect 493910 633980 494530 633985
rect 493910 633360 493920 633980
rect 494520 633360 494530 633980
rect 493910 633355 494530 633360
rect 570200 631000 572000 643000
rect 580000 631000 582858 643000
rect 570200 629814 582858 631000
rect 570200 629800 582262 629814
rect 427731 627183 427741 629635
rect 439681 628990 439691 629635
rect 439681 627828 492245 628990
rect 439681 627183 439691 627828
rect 490970 626707 491712 626722
rect 490970 626643 490990 626707
rect 491054 626694 491712 626707
rect 491054 626689 491728 626694
rect 491054 626643 491662 626689
rect 490970 626633 491662 626643
rect 491718 626633 491728 626689
rect 490970 626628 491728 626633
rect 490970 626622 491712 626628
rect 490968 626545 491722 626550
rect 490968 626531 491656 626545
rect 490968 626467 490992 626531
rect 491056 626489 491656 626531
rect 491712 626489 491722 626545
rect 491056 626484 491722 626489
rect 491056 626467 491710 626484
rect 490968 626450 491710 626467
rect 291988 595121 487458 595469
rect 291988 594419 486464 595121
rect 487165 594419 487458 595121
rect 291988 594152 487458 594419
rect 443868 592894 445765 592903
rect 294628 592621 446728 592894
rect 294628 591743 443717 592621
rect 446222 591743 446728 592621
rect 294628 591488 446728 591743
rect 294628 591472 443702 591488
rect 446425 591472 446728 591488
rect 490416 586522 490426 589002
rect 490676 586522 490686 589002
rect 581138 587168 581148 587930
rect 581394 587928 581404 587930
rect 581394 587168 582714 587928
rect 523864 569681 523874 569950
rect 515889 569669 523874 569681
rect 515889 569455 515905 569669
rect 516059 569455 523874 569669
rect 515889 569442 523874 569455
rect 523864 569133 523874 569442
rect 527538 569133 527548 569950
rect 413308 566115 413318 567480
rect 417373 566607 417383 567480
rect 443868 566607 445765 566635
rect 417373 566596 491700 566607
rect 417373 566115 491505 566596
rect 417083 565941 491505 566115
rect 417083 565910 443148 565941
rect 446540 565936 491505 565941
rect 491689 565936 491700 566596
rect 446540 565910 491700 565936
rect 486181 559030 487344 559035
rect 486181 557812 486191 559030
rect 487334 558751 487344 559030
rect 495615 558751 495733 560106
rect 536894 559292 536904 559337
rect 513760 559279 536904 559292
rect 513760 559215 513778 559279
rect 513842 559233 536904 559279
rect 537239 559233 537249 559337
rect 513842 559215 537229 559233
rect 513760 559204 537229 559215
rect 547500 559142 547510 559184
rect 496792 559132 547510 559142
rect 496792 559068 496813 559132
rect 496877 559068 547510 559132
rect 496792 559054 547510 559068
rect 547500 559028 547510 559054
rect 547652 559028 547662 559184
rect 487334 557932 495741 558751
rect 487334 557812 487344 557932
rect 486181 557807 487344 557812
rect 401584 467823 403762 468039
rect 400108 466110 400118 467823
rect 401862 466110 403762 467823
rect 401584 413613 403762 466110
rect 443872 455747 445769 456513
rect 443750 455126 443760 455747
rect 445837 455126 445847 455747
rect 443872 453650 445769 455126
rect 443868 453628 445769 453650
rect 443868 450765 445765 453628
rect 446134 453584 461586 453589
rect 446134 451623 446144 453584
rect 461576 451623 461586 453584
rect 446134 451618 461586 451623
rect 443868 450566 444699 450765
rect 445166 450566 445765 450765
rect 443868 450532 445765 450566
rect 426670 449375 426680 450393
rect 440871 449885 440881 450393
rect 440871 449531 443842 449885
rect 440871 449526 443844 449531
rect 440871 449375 440881 449526
rect 443649 449514 443844 449526
rect 443649 418942 443847 449514
rect 401582 412519 403764 413613
rect 401582 412425 403648 412519
rect 403740 412425 403764 412519
rect 401582 412398 403764 412425
rect 401669 411980 403841 412237
rect 401669 411886 403659 411980
rect 403751 411886 403841 411980
rect 401669 361852 403841 411886
rect 441966 382352 441976 386778
rect 442336 382352 442346 386778
rect 400136 360139 400146 361852
rect 401890 360139 403841 361852
rect 401669 360023 403841 360139
rect 473797 355440 473807 355592
rect 467461 355425 473807 355440
rect 467461 355277 467471 355425
rect 467538 355277 473807 355425
rect 467461 355271 473807 355277
rect 477651 355271 477661 355592
rect 467461 355269 474072 355271
rect 413248 351802 413258 352663
rect 418042 352485 418052 352663
rect 418042 352478 443261 352485
rect 418042 352473 443264 352478
rect 418042 352045 443150 352473
rect 443254 352045 443264 352473
rect 418042 352040 443264 352045
rect 418042 352030 443261 352040
rect 418042 351802 418052 352030
rect 535689 345624 535699 345920
rect 473196 345598 535699 345624
rect 473196 345534 473216 345598
rect 473280 345534 535699 345598
rect 473196 345519 535699 345534
rect 535689 345427 535699 345519
rect 540805 345427 540815 345920
rect 491824 344559 535221 344560
rect 546047 344559 546057 344834
rect 448355 344544 546057 344559
rect 448355 344480 448374 344544
rect 448438 344480 546057 344544
rect 448355 344466 546057 344480
rect 448355 344465 535221 344466
rect 448355 344464 491835 344465
rect 546047 344326 546057 344466
rect 551617 344326 551627 344834
<< via3 >>
rect 474059 700807 477386 702380
rect 511000 694000 525000 702000
rect 537573 699875 540501 702106
rect 548589 678122 551656 681190
rect 493920 633360 494520 633980
rect 572000 631000 580000 643000
rect 427741 627183 439681 629635
rect 490990 626643 491054 626707
rect 490992 626467 491056 626531
rect 443717 591743 446222 592621
rect 490426 586522 490676 589002
rect 581148 587168 581394 587930
rect 523874 569133 527538 569950
rect 413318 566115 417373 567480
rect 536904 559233 537239 559337
rect 547510 559028 547652 559184
rect 400118 466110 401862 467823
rect 443760 455126 445837 455747
rect 446144 451623 461576 453584
rect 426680 449375 440871 450393
rect 441976 382352 442336 386778
rect 400146 360139 401890 361852
rect 473807 355271 477651 355592
rect 413258 351802 418042 352663
rect 535699 345427 540805 345920
rect 546057 344326 551617 344834
<< metal4 >>
rect 216408 701118 233422 703354
rect 318686 702196 335618 702676
rect 216456 624926 233394 701118
rect 318718 628567 335656 702196
rect 412976 702036 418408 702596
rect 473692 702380 477800 702424
rect 473692 702320 474059 702380
rect 318718 626984 319826 628567
rect 334706 626984 335656 628567
rect 318718 625718 335656 626984
rect 216456 622868 217881 624926
rect 232603 622868 233394 624926
rect 216456 621602 233394 622868
rect 412985 567480 418341 702036
rect 473693 700807 474059 702320
rect 477386 700807 477803 702380
rect 510002 702246 525998 702538
rect 426493 691654 441057 693607
rect 426493 691459 428802 691654
rect 426490 679221 428802 691459
rect 439991 679221 441057 691654
rect 412985 566115 413318 567480
rect 417373 566115 418341 567480
rect 400117 467823 401863 467824
rect 400117 466110 400118 467823
rect 401862 466110 401863 467823
rect 400117 466109 401863 466110
rect 400145 361852 401891 361853
rect 400145 360139 400146 361852
rect 401890 360139 401891 361852
rect 400145 360138 401891 360139
rect 412985 359017 418341 566115
rect 419918 664392 424966 665528
rect 419918 659652 420524 664392
rect 424428 659652 424966 664392
rect 419918 418550 424966 659652
rect 426490 629635 441057 679221
rect 473693 657000 477803 700807
rect 510000 702173 526000 702246
rect 510000 702000 511182 702173
rect 510000 694000 511000 702000
rect 510000 689303 511182 694000
rect 525301 689303 526000 702173
rect 510000 683200 526000 689303
rect 536032 702106 541241 702380
rect 536032 699875 537573 702106
rect 540501 699875 541241 702106
rect 473693 649762 474474 657000
rect 477728 649762 477803 657000
rect 426490 627183 427741 629635
rect 439681 627183 441057 629635
rect 426490 451355 441057 627183
rect 448886 645202 464003 646531
rect 448886 631579 451046 645202
rect 463339 631579 464003 645202
rect 443481 592621 446243 592793
rect 443481 591743 443717 592621
rect 446222 591743 446243 592621
rect 443481 455747 446243 591743
rect 443481 455126 443760 455747
rect 445837 455126 446243 455747
rect 443481 454827 446243 455126
rect 448886 453585 464003 631579
rect 446143 453584 464003 453585
rect 446143 451623 446144 453584
rect 461576 451623 464003 453584
rect 446143 451622 464003 451623
rect 426490 450393 441054 451355
rect 448886 451335 464003 451622
rect 426490 449375 426680 450393
rect 440871 449375 441054 450393
rect 426490 449207 441054 449375
rect 419918 418232 420512 418550
rect 424392 418232 424966 418550
rect 419918 417788 424966 418232
rect 441975 386778 442337 386779
rect 441975 382352 441976 386778
rect 442336 382352 442337 386778
rect 441975 382351 442337 382352
rect 412954 357954 418341 359017
rect 412954 352663 418320 357954
rect 473693 355592 477803 649762
rect 493072 632978 493142 658010
rect 523682 655766 527778 656215
rect 523682 650604 524748 655766
rect 527329 650604 527778 655766
rect 493919 633980 494521 633981
rect 493919 633360 493920 633980
rect 494520 633360 494521 633980
rect 493919 633359 494521 633360
rect 490977 626707 491090 627229
rect 490977 626643 490990 626707
rect 491054 626643 491090 626707
rect 490977 626630 491090 626643
rect 490912 626532 491055 626547
rect 490912 626531 491057 626532
rect 490912 626467 490992 626531
rect 491056 626467 491057 626531
rect 490912 626466 491057 626467
rect 490912 624574 491055 626466
rect 490999 624549 491055 624574
rect 490999 624338 491057 624549
rect 490425 589002 490677 589003
rect 490425 586522 490426 589002
rect 490676 586522 490677 589002
rect 490425 586521 490677 586522
rect 523682 569950 527778 650604
rect 523682 569133 523874 569950
rect 527538 569133 527778 569950
rect 523682 566832 527778 569133
rect 536032 562758 541241 699875
rect 473693 355271 473807 355592
rect 477651 355271 477803 355592
rect 473693 355203 477803 355271
rect 535604 559337 541241 562758
rect 545992 681190 551755 682997
rect 545992 678122 548589 681190
rect 551656 678122 551755 681190
rect 545992 562330 551755 678122
rect 570000 643000 582000 645000
rect 570000 631000 572000 643000
rect 580000 631000 582000 643000
rect 570000 630000 582000 631000
rect 535604 559233 536904 559337
rect 537239 559248 541241 559337
rect 537239 559233 540970 559248
rect 412954 351802 413258 352663
rect 418042 351802 418320 352663
rect 412954 351473 418320 351802
rect 535604 347330 540970 559233
rect 545948 559184 551755 562330
rect 545948 559028 547510 559184
rect 547652 559028 551755 559184
rect 545948 558353 551755 559028
rect 560006 588286 564916 589148
rect 560006 587038 561644 588286
rect 563946 587038 564916 588286
rect 581147 587930 581395 587931
rect 581147 587168 581148 587930
rect 581394 587168 581395 587930
rect 581147 587167 581395 587168
rect 535604 346960 540973 347330
rect 535605 345920 540973 346960
rect 535605 345427 535699 345920
rect 540805 345427 540973 345920
rect 535605 345350 540973 345427
rect 545948 344834 551744 558353
rect 560006 386392 564916 587038
rect 560006 382888 560754 386392
rect 563860 382888 564916 386392
rect 560006 382170 564916 382888
rect 545948 344326 546057 344834
rect 551617 344326 551744 344834
rect 545948 342093 551744 344326
<< via4 >>
rect 319826 626984 334706 628567
rect 217881 622868 232603 624926
rect 428802 679221 439991 691654
rect 400118 466110 401862 467823
rect 400146 360139 401890 361852
rect 420524 659652 424428 664392
rect 511182 702000 525301 702173
rect 511182 694000 525000 702000
rect 525000 694000 525301 702000
rect 511182 689303 525301 694000
rect 492836 658010 493638 666470
rect 474474 649762 477728 657000
rect 451046 631579 463339 645202
rect 420512 418232 424392 418550
rect 444600 418384 444836 418620
rect 441976 382352 442336 386778
rect 524748 650604 527329 655766
rect 493920 633360 494520 633980
rect 490940 627229 491176 627465
rect 490763 624338 490999 624574
rect 490426 586522 490676 589002
rect 572000 631000 580000 643000
rect 561644 587038 563946 588286
rect 581148 587168 581394 587930
rect 560754 382888 563860 386392
<< metal5 >>
rect 511158 702173 525325 702197
rect 511158 694673 511182 702173
rect 426493 691654 511182 694673
rect 426493 679221 428802 691654
rect 439991 689303 511182 691654
rect 525301 694673 525325 702173
rect 525301 689303 525419 694673
rect 439991 679221 525419 689303
rect 426493 677090 525419 679221
rect 165400 666470 498120 666708
rect 165400 664392 492836 666470
rect 165400 659652 420524 664392
rect 424428 659652 492836 664392
rect 165400 658010 492836 659652
rect 493638 658010 498120 666470
rect 165400 657886 498120 658010
rect 474450 657000 477752 657024
rect 474450 649762 474474 657000
rect 477728 656197 477752 657000
rect 477728 655766 527767 656197
rect 477728 650604 524748 655766
rect 527329 650604 527767 655766
rect 477728 650182 527767 650604
rect 477728 649762 477752 650182
rect 474450 649738 477752 649762
rect 449052 646960 526532 647014
rect 560200 646960 582000 647000
rect 449052 645202 582000 646960
rect 449052 631579 451046 645202
rect 463339 643000 582000 645202
rect 463339 633980 572000 643000
rect 463339 633360 493920 633980
rect 494520 633360 572000 633980
rect 463339 631579 572000 633360
rect 449052 631000 572000 631579
rect 580000 631000 582000 643000
rect 449052 630084 582000 631000
rect 485200 630030 582000 630084
rect 560200 630000 582000 630030
rect 331386 628591 491233 628693
rect 319802 628567 491233 628591
rect 319802 626984 319826 628567
rect 334706 627465 491233 628567
rect 334706 627229 490940 627465
rect 491176 627229 491233 627465
rect 334706 627195 491233 627229
rect 334706 626984 334730 627195
rect 319802 626960 334730 626984
rect 217857 624926 232627 624950
rect 217857 622868 217881 624926
rect 232603 624611 232627 624926
rect 232603 624574 491025 624611
rect 232603 624338 490763 624574
rect 490999 624338 491025 624574
rect 232603 622964 491025 624338
rect 232603 622868 232627 622964
rect 217857 622844 232627 622868
rect 489376 589002 581822 589152
rect 489376 586522 490426 589002
rect 490676 588286 581822 589002
rect 490676 587038 561644 588286
rect 563946 587930 581822 588286
rect 563946 587168 581148 587930
rect 581394 587168 581822 587930
rect 563946 587038 581822 587168
rect 490676 586522 581822 587038
rect 489376 586448 581822 586522
rect 400094 467823 401886 467847
rect 400094 466110 400118 467823
rect 401862 466110 401886 467823
rect 400094 466086 401886 466110
rect 423776 418620 444862 418654
rect 423776 418574 444600 418620
rect 420488 418550 444600 418574
rect 420488 418232 420512 418550
rect 424392 418384 444600 418550
rect 444836 418384 444862 418620
rect 424392 418266 444862 418384
rect 424392 418232 424416 418266
rect 420488 418208 424416 418232
rect 441342 386778 564420 386914
rect 441342 382352 441976 386778
rect 442336 386392 564420 386778
rect 442336 382888 560754 386392
rect 563860 382888 564420 386392
rect 442336 382352 564420 382888
rect 441342 382166 564420 382352
rect 399700 361852 401998 362010
rect 399700 360139 400146 361852
rect 401890 360139 401998 361852
rect 399700 360009 401998 360139
<< comment >>
rect 584000 323622 584100 350000
use top  top_0
timestamp 1662990520
transform 1 0 443353 0 1 404933
box -2734 -60442 26330 14173
use top  top_1
timestamp 1662990520
transform 1 0 491794 0 1 619522
box -2734 -60442 26330 14173
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
