magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -346 1454 1506 1586
rect -346 206 -214 1454
rect 1374 206 1506 1454
rect -346 74 1506 206
rect -346 -1174 -214 74
rect 1374 -1174 1506 74
rect -346 -1306 1506 -1174
<< psubdiff >>
rect -320 1537 1480 1560
rect -320 1503 -195 1537
rect -161 1503 -127 1537
rect -93 1503 -59 1537
rect -25 1503 265 1537
rect 299 1503 333 1537
rect 367 1503 401 1537
rect 435 1503 725 1537
rect 759 1503 793 1537
rect 827 1503 861 1537
rect 895 1503 1185 1537
rect 1219 1503 1253 1537
rect 1287 1503 1321 1537
rect 1355 1503 1480 1537
rect -320 1480 1480 1503
rect -320 1175 -240 1480
rect -320 1141 -297 1175
rect -263 1141 -240 1175
rect -320 1107 -240 1141
rect -320 1073 -297 1107
rect -263 1073 -240 1107
rect -320 1039 -240 1073
rect -320 1005 -297 1039
rect -263 1005 -240 1039
rect -320 695 -240 1005
rect -320 661 -297 695
rect -263 661 -240 695
rect -320 627 -240 661
rect -320 593 -297 627
rect -263 593 -240 627
rect -320 559 -240 593
rect -320 525 -297 559
rect -263 525 -240 559
rect -320 180 -240 525
rect 1400 1175 1480 1480
rect 1400 1141 1423 1175
rect 1457 1141 1480 1175
rect 1400 1107 1480 1141
rect 1400 1073 1423 1107
rect 1457 1073 1480 1107
rect 1400 1039 1480 1073
rect 1400 1005 1423 1039
rect 1457 1005 1480 1039
rect 1400 695 1480 1005
rect 1400 661 1423 695
rect 1457 661 1480 695
rect 1400 627 1480 661
rect 1400 593 1423 627
rect 1457 593 1480 627
rect 1400 559 1480 593
rect 1400 525 1423 559
rect 1457 525 1480 559
rect 1400 180 1480 525
rect -320 157 1480 180
rect -320 123 -195 157
rect -161 123 -127 157
rect -93 123 -59 157
rect -25 123 265 157
rect 299 123 333 157
rect 367 123 401 157
rect 435 123 725 157
rect 759 123 793 157
rect 827 123 861 157
rect 895 123 1185 157
rect 1219 123 1253 157
rect 1287 123 1321 157
rect 1355 123 1480 157
rect -320 100 1480 123
rect -320 -165 -240 100
rect -320 -199 -297 -165
rect -263 -199 -240 -165
rect -320 -233 -240 -199
rect -320 -267 -297 -233
rect -263 -267 -240 -233
rect -320 -301 -240 -267
rect -320 -335 -297 -301
rect -263 -335 -240 -301
rect -320 -725 -240 -335
rect -320 -759 -297 -725
rect -263 -759 -240 -725
rect -320 -793 -240 -759
rect -320 -827 -297 -793
rect -263 -827 -240 -793
rect -320 -861 -240 -827
rect -320 -895 -297 -861
rect -263 -895 -240 -861
rect -320 -1200 -240 -895
rect 1400 -165 1480 100
rect 1400 -199 1423 -165
rect 1457 -199 1480 -165
rect 1400 -233 1480 -199
rect 1400 -267 1423 -233
rect 1457 -267 1480 -233
rect 1400 -301 1480 -267
rect 1400 -335 1423 -301
rect 1457 -335 1480 -301
rect 1400 -725 1480 -335
rect 1400 -759 1423 -725
rect 1457 -759 1480 -725
rect 1400 -793 1480 -759
rect 1400 -827 1423 -793
rect 1457 -827 1480 -793
rect 1400 -861 1480 -827
rect 1400 -895 1423 -861
rect 1457 -895 1480 -861
rect 1400 -1200 1480 -895
rect -320 -1223 1480 -1200
rect -320 -1257 -195 -1223
rect -161 -1257 -127 -1223
rect -93 -1257 -59 -1223
rect -25 -1257 265 -1223
rect 299 -1257 333 -1223
rect 367 -1257 401 -1223
rect 435 -1257 725 -1223
rect 759 -1257 793 -1223
rect 827 -1257 861 -1223
rect 895 -1257 1185 -1223
rect 1219 -1257 1253 -1223
rect 1287 -1257 1321 -1223
rect 1355 -1257 1480 -1223
rect -320 -1280 1480 -1257
<< psubdiffcont >>
rect -195 1503 -161 1537
rect -127 1503 -93 1537
rect -59 1503 -25 1537
rect 265 1503 299 1537
rect 333 1503 367 1537
rect 401 1503 435 1537
rect 725 1503 759 1537
rect 793 1503 827 1537
rect 861 1503 895 1537
rect 1185 1503 1219 1537
rect 1253 1503 1287 1537
rect 1321 1503 1355 1537
rect -297 1141 -263 1175
rect -297 1073 -263 1107
rect -297 1005 -263 1039
rect -297 661 -263 695
rect -297 593 -263 627
rect -297 525 -263 559
rect 1423 1141 1457 1175
rect 1423 1073 1457 1107
rect 1423 1005 1457 1039
rect 1423 661 1457 695
rect 1423 593 1457 627
rect 1423 525 1457 559
rect -195 123 -161 157
rect -127 123 -93 157
rect -59 123 -25 157
rect 265 123 299 157
rect 333 123 367 157
rect 401 123 435 157
rect 725 123 759 157
rect 793 123 827 157
rect 861 123 895 157
rect 1185 123 1219 157
rect 1253 123 1287 157
rect 1321 123 1355 157
rect -297 -199 -263 -165
rect -297 -267 -263 -233
rect -297 -335 -263 -301
rect -297 -759 -263 -725
rect -297 -827 -263 -793
rect -297 -895 -263 -861
rect 1423 -199 1457 -165
rect 1423 -267 1457 -233
rect 1423 -335 1457 -301
rect 1423 -759 1457 -725
rect 1423 -827 1457 -793
rect 1423 -895 1457 -861
rect -195 -1257 -161 -1223
rect -127 -1257 -93 -1223
rect -59 -1257 -25 -1223
rect 265 -1257 299 -1223
rect 333 -1257 367 -1223
rect 401 -1257 435 -1223
rect 725 -1257 759 -1223
rect 793 -1257 827 -1223
rect 861 -1257 895 -1223
rect 1185 -1257 1219 -1223
rect 1253 -1257 1287 -1223
rect 1321 -1257 1355 -1223
<< locali >>
rect -320 1537 1480 1560
rect -320 1503 -199 1537
rect -161 1503 -127 1537
rect -93 1503 -59 1537
rect -21 1503 261 1537
rect 299 1503 333 1537
rect 367 1503 401 1537
rect 439 1503 721 1537
rect 759 1503 793 1537
rect 827 1503 861 1537
rect 899 1503 1181 1537
rect 1219 1503 1253 1537
rect 1287 1503 1321 1537
rect 1359 1503 1480 1537
rect -320 1480 1480 1503
rect -320 1179 -240 1480
rect -320 1141 -297 1179
rect -263 1141 -240 1179
rect -320 1107 -240 1141
rect -320 1073 -297 1107
rect -263 1073 -240 1107
rect -320 1039 -240 1073
rect -320 1001 -297 1039
rect -263 1001 -240 1039
rect -320 699 -240 1001
rect -320 661 -297 699
rect -263 661 -240 699
rect -320 627 -240 661
rect -320 593 -297 627
rect -263 593 -240 627
rect -320 559 -240 593
rect -320 521 -297 559
rect -263 521 -240 559
rect -320 180 -240 521
rect 1400 1179 1480 1480
rect 1400 1141 1423 1179
rect 1457 1141 1480 1179
rect 1400 1107 1480 1141
rect 1400 1073 1423 1107
rect 1457 1073 1480 1107
rect 1400 1039 1480 1073
rect 1400 1001 1423 1039
rect 1457 1001 1480 1039
rect 1400 699 1480 1001
rect 1400 661 1423 699
rect 1457 661 1480 699
rect 1400 627 1480 661
rect 1400 593 1423 627
rect 1457 593 1480 627
rect 1400 559 1480 593
rect 1400 521 1423 559
rect 1457 521 1480 559
rect 1400 180 1480 521
rect -320 157 1480 180
rect -320 123 -195 157
rect -161 123 -127 157
rect -93 123 -59 157
rect -25 123 265 157
rect 299 123 333 157
rect 367 123 401 157
rect 435 123 725 157
rect 759 123 793 157
rect 827 123 861 157
rect 895 123 1185 157
rect 1219 123 1253 157
rect 1287 123 1321 157
rect 1355 123 1480 157
rect -320 100 1480 123
rect -320 -161 -240 100
rect -320 -199 -297 -161
rect -263 -199 -240 -161
rect -320 -233 -240 -199
rect -320 -267 -297 -233
rect -263 -267 -240 -233
rect -320 -301 -240 -267
rect -320 -339 -297 -301
rect -263 -339 -240 -301
rect -320 -721 -240 -339
rect -320 -759 -297 -721
rect -263 -759 -240 -721
rect -320 -793 -240 -759
rect -320 -827 -297 -793
rect -263 -827 -240 -793
rect -320 -861 -240 -827
rect -320 -899 -297 -861
rect -263 -899 -240 -861
rect -320 -1200 -240 -899
rect 1400 -161 1480 100
rect 1400 -199 1423 -161
rect 1457 -199 1480 -161
rect 1400 -233 1480 -199
rect 1400 -267 1423 -233
rect 1457 -267 1480 -233
rect 1400 -301 1480 -267
rect 1400 -339 1423 -301
rect 1457 -339 1480 -301
rect 1400 -721 1480 -339
rect 1400 -759 1423 -721
rect 1457 -759 1480 -721
rect 1400 -793 1480 -759
rect 1400 -827 1423 -793
rect 1457 -827 1480 -793
rect 1400 -861 1480 -827
rect 1400 -899 1423 -861
rect 1457 -899 1480 -861
rect 1400 -1200 1480 -899
rect -320 -1223 1480 -1200
rect -320 -1257 -199 -1223
rect -161 -1257 -127 -1223
rect -93 -1257 -59 -1223
rect -21 -1257 261 -1223
rect 299 -1257 333 -1223
rect 367 -1257 401 -1223
rect 439 -1257 721 -1223
rect 759 -1257 793 -1223
rect 827 -1257 861 -1223
rect 899 -1257 1181 -1223
rect 1219 -1257 1253 -1223
rect 1287 -1257 1321 -1223
rect 1359 -1257 1480 -1223
rect -320 -1280 1480 -1257
<< viali >>
rect -199 1503 -195 1537
rect -195 1503 -165 1537
rect -127 1503 -93 1537
rect -55 1503 -25 1537
rect -25 1503 -21 1537
rect 261 1503 265 1537
rect 265 1503 295 1537
rect 333 1503 367 1537
rect 405 1503 435 1537
rect 435 1503 439 1537
rect 721 1503 725 1537
rect 725 1503 755 1537
rect 793 1503 827 1537
rect 865 1503 895 1537
rect 895 1503 899 1537
rect 1181 1503 1185 1537
rect 1185 1503 1215 1537
rect 1253 1503 1287 1537
rect 1325 1503 1355 1537
rect 1355 1503 1359 1537
rect -297 1175 -263 1179
rect -297 1145 -263 1175
rect -297 1073 -263 1107
rect -297 1005 -263 1035
rect -297 1001 -263 1005
rect -297 695 -263 699
rect -297 665 -263 695
rect -297 593 -263 627
rect -297 525 -263 555
rect -297 521 -263 525
rect 1423 1175 1457 1179
rect 1423 1145 1457 1175
rect 1423 1073 1457 1107
rect 1423 1005 1457 1035
rect 1423 1001 1457 1005
rect 1423 695 1457 699
rect 1423 665 1457 695
rect 1423 593 1457 627
rect 1423 525 1457 555
rect 1423 521 1457 525
rect -297 -165 -263 -161
rect -297 -195 -263 -165
rect -297 -267 -263 -233
rect -297 -335 -263 -305
rect -297 -339 -263 -335
rect -297 -725 -263 -721
rect -297 -755 -263 -725
rect -297 -827 -263 -793
rect -297 -895 -263 -865
rect -297 -899 -263 -895
rect 1423 -165 1457 -161
rect 1423 -195 1457 -165
rect 1423 -267 1457 -233
rect 1423 -335 1457 -305
rect 1423 -339 1457 -335
rect 1423 -725 1457 -721
rect 1423 -755 1457 -725
rect 1423 -827 1457 -793
rect 1423 -895 1457 -865
rect 1423 -899 1457 -895
rect -199 -1257 -195 -1223
rect -195 -1257 -165 -1223
rect -127 -1257 -93 -1223
rect -55 -1257 -25 -1223
rect -25 -1257 -21 -1223
rect 261 -1257 265 -1223
rect 265 -1257 295 -1223
rect 333 -1257 367 -1223
rect 405 -1257 435 -1223
rect 435 -1257 439 -1223
rect 721 -1257 725 -1223
rect 725 -1257 755 -1223
rect 793 -1257 827 -1223
rect 865 -1257 895 -1223
rect 895 -1257 899 -1223
rect 1181 -1257 1185 -1223
rect 1185 -1257 1215 -1223
rect 1253 -1257 1287 -1223
rect 1325 -1257 1355 -1223
rect 1355 -1257 1359 -1223
<< metal1 >>
rect -320 1537 1480 1560
rect -320 1503 -199 1537
rect -165 1503 -127 1537
rect -93 1503 -55 1537
rect -21 1503 261 1537
rect 295 1503 333 1537
rect 367 1503 405 1537
rect 439 1503 721 1537
rect 755 1503 793 1537
rect 827 1503 865 1537
rect 899 1503 1181 1537
rect 1215 1503 1253 1537
rect 1287 1503 1325 1537
rect 1359 1503 1480 1537
rect -320 1480 1480 1503
rect -320 1179 -240 1480
rect 30 1336 110 1340
rect 30 1284 44 1336
rect 96 1284 110 1336
rect 30 1280 110 1284
rect 1060 1336 1140 1340
rect 1060 1284 1074 1336
rect 1126 1284 1140 1336
rect 1060 1280 1140 1284
rect -320 1145 -297 1179
rect -263 1145 -240 1179
rect -320 1107 -240 1145
rect -320 1073 -297 1107
rect -263 1073 -240 1107
rect -320 1035 -240 1073
rect -320 1001 -297 1035
rect -263 1001 -240 1035
rect -320 699 -240 1001
rect 1400 1179 1480 1480
rect 1400 1145 1423 1179
rect 1457 1145 1480 1179
rect 1400 1107 1480 1145
rect 1400 1073 1423 1107
rect 1457 1073 1480 1107
rect 1400 1035 1480 1073
rect 1400 1001 1423 1035
rect 1457 1001 1480 1035
rect 280 896 370 910
rect 280 844 299 896
rect 351 844 370 896
rect 280 830 370 844
rect 790 896 880 910
rect 790 844 809 896
rect 861 844 880 896
rect 790 830 880 844
rect -320 665 -297 699
rect -263 665 -240 699
rect -320 627 -240 665
rect -320 593 -297 627
rect -263 593 -240 627
rect -320 555 -240 593
rect -320 521 -297 555
rect -263 521 -240 555
rect -320 -161 -240 521
rect 1400 699 1480 1001
rect 1400 665 1423 699
rect 1457 665 1480 699
rect 1400 627 1480 665
rect 1400 593 1423 627
rect 1457 593 1480 627
rect 1400 555 1480 593
rect 1400 521 1423 555
rect 1457 521 1480 555
rect 544 494 624 498
rect 544 442 558 494
rect 610 442 624 494
rect 544 438 624 442
rect 160 256 240 400
rect 160 204 174 256
rect 226 204 240 256
rect 160 200 240 204
rect 160 76 240 80
rect 160 24 174 76
rect 226 24 240 76
rect 160 -120 240 24
rect 430 76 510 400
rect 551 360 619 406
rect 430 24 444 76
rect 496 24 510 76
rect 430 20 510 24
rect 660 256 740 260
rect 660 204 674 256
rect 726 204 740 256
rect 551 -122 619 -76
rect 660 -120 740 204
rect 930 256 1010 400
rect 930 204 944 256
rect 996 204 1010 256
rect 930 200 1010 204
rect 930 76 1010 80
rect 930 24 944 76
rect 996 24 1010 76
rect 930 -120 1010 24
rect -320 -195 -297 -161
rect -263 -195 -240 -161
rect -320 -233 -240 -195
rect 545 -158 625 -154
rect 545 -210 559 -158
rect 611 -210 625 -158
rect 545 -214 625 -210
rect 1400 -161 1480 521
rect 1400 -195 1423 -161
rect 1457 -195 1480 -161
rect -320 -267 -297 -233
rect -263 -267 -240 -233
rect -320 -305 -240 -267
rect -320 -339 -297 -305
rect -263 -339 -240 -305
rect -320 -721 -240 -339
rect 1400 -233 1480 -195
rect 1400 -267 1423 -233
rect 1457 -267 1480 -233
rect 1400 -305 1480 -267
rect 1400 -339 1423 -305
rect 1457 -339 1480 -305
rect 280 -604 370 -590
rect 280 -656 299 -604
rect 351 -656 370 -604
rect 280 -670 370 -656
rect 790 -604 880 -590
rect 790 -656 809 -604
rect 861 -656 880 -604
rect 790 -670 880 -656
rect -320 -755 -297 -721
rect -263 -755 -240 -721
rect -320 -793 -240 -755
rect -320 -827 -297 -793
rect -263 -827 -240 -793
rect -320 -865 -240 -827
rect -320 -899 -297 -865
rect -263 -899 -240 -865
rect -320 -1200 -240 -899
rect 1400 -721 1480 -339
rect 1400 -755 1423 -721
rect 1457 -755 1480 -721
rect 1400 -793 1480 -755
rect 1400 -827 1423 -793
rect 1457 -827 1480 -793
rect 1400 -865 1480 -827
rect 1400 -899 1423 -865
rect 1457 -899 1480 -865
rect 30 -1004 110 -1000
rect 30 -1056 44 -1004
rect 96 -1056 110 -1004
rect 30 -1060 110 -1056
rect 1060 -1004 1140 -1000
rect 1060 -1056 1074 -1004
rect 1126 -1056 1140 -1004
rect 1060 -1060 1140 -1056
rect 1400 -1200 1480 -899
rect -320 -1223 1480 -1200
rect -320 -1257 -199 -1223
rect -165 -1257 -127 -1223
rect -93 -1257 -55 -1223
rect -21 -1257 261 -1223
rect 295 -1257 333 -1223
rect 367 -1257 405 -1223
rect 439 -1257 721 -1223
rect 755 -1257 793 -1223
rect 827 -1257 865 -1223
rect 899 -1257 1181 -1223
rect 1215 -1257 1253 -1223
rect 1287 -1257 1325 -1223
rect 1359 -1257 1480 -1223
rect -320 -1280 1480 -1257
<< via1 >>
rect 44 1284 96 1336
rect 1074 1284 1126 1336
rect 299 844 351 896
rect 809 844 861 896
rect 558 442 610 494
rect 174 204 226 256
rect 174 24 226 76
rect 444 24 496 76
rect 674 204 726 256
rect 944 204 996 256
rect 944 24 996 76
rect 559 -210 611 -158
rect 299 -656 351 -604
rect 809 -656 861 -604
rect 44 -1056 96 -1004
rect 1074 -1056 1126 -1004
<< metal2 >>
rect 40 1336 1266 1350
rect 40 1284 44 1336
rect 96 1284 1074 1336
rect 1126 1284 1266 1336
rect 40 1270 1266 1284
rect 290 898 870 920
rect 290 842 297 898
rect 353 896 870 898
rect 353 844 809 896
rect 861 844 870 896
rect 353 842 870 844
rect 290 820 870 842
rect -98 494 614 508
rect -98 442 558 494
rect 610 442 614 494
rect -98 428 614 442
rect -98 -990 -30 428
rect 170 256 1000 270
rect 170 204 174 256
rect 226 204 674 256
rect 726 204 944 256
rect 996 204 1000 256
rect 170 190 1000 204
rect 170 76 1000 90
rect 170 24 174 76
rect 226 24 444 76
rect 496 24 944 76
rect 996 24 1000 76
rect 170 10 1000 24
rect 1198 -144 1266 1270
rect 554 -158 1266 -144
rect 554 -210 559 -158
rect 611 -210 1266 -158
rect 554 -224 1266 -210
rect 290 -602 870 -580
rect 290 -658 297 -602
rect 353 -604 870 -602
rect 353 -656 809 -604
rect 861 -656 870 -604
rect 353 -658 870 -656
rect 290 -680 870 -658
rect -98 -1004 1130 -990
rect -98 -1056 44 -1004
rect 96 -1056 1074 -1004
rect 1126 -1056 1130 -1004
rect -98 -1070 1130 -1056
<< via2 >>
rect 297 896 353 898
rect 297 844 299 896
rect 299 844 351 896
rect 351 844 353 896
rect 297 842 353 844
rect 297 -604 353 -602
rect 297 -656 299 -604
rect 299 -656 351 -604
rect 351 -656 353 -604
rect 297 -658 353 -656
<< metal3 >>
rect 280 898 380 920
rect 280 842 297 898
rect 353 842 380 898
rect 280 180 380 842
rect -360 100 380 180
rect 280 -602 380 100
rect 280 -658 297 -602
rect 353 -658 380 -602
rect 280 -680 380 -658
use sky130_fd_pr__nfet_01v8_lvt_A5VCMN  sky130_fd_pr__nfet_01v8_lvt_A5VCMN_0
timestamp 1663011646
transform 1 0 585 0 1 -573
box -571 -507 571 507
use sky130_fd_pr__nfet_01v8_lvt_E96B6C  sky130_fd_pr__nfet_01v8_lvt_E96B6C_0
timestamp 1663011646
transform 1 0 585 0 1 857
box -571 -507 571 507
<< end >>
