magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal1 >>
rect 522 3002 622 3026
rect 522 2950 546 3002
rect 598 2950 622 3002
rect 522 2926 622 2950
rect 1438 3002 1538 3026
rect 1438 2950 1462 3002
rect 1514 2950 1538 3002
rect 1438 2926 1538 2950
rect 2352 3002 2452 3026
rect 2352 2950 2376 3002
rect 2428 2950 2452 3002
rect 2352 2926 2452 2950
rect 1465 2916 1471 2926
rect 1505 2916 1511 2926
rect 2379 2916 2385 2926
rect 2419 2916 2425 2926
rect 1921 2536 1927 2546
rect 1961 2536 1967 2546
rect 1007 2524 1013 2534
rect 1047 2524 1053 2534
rect 64 2500 164 2524
rect 64 2448 88 2500
rect 140 2448 164 2500
rect 64 2424 164 2448
rect 980 2500 1080 2524
rect 980 2448 1004 2500
rect 1056 2448 1080 2500
rect 980 2424 1080 2448
rect 1894 2512 1994 2536
rect 1894 2460 1918 2512
rect 1970 2460 1994 2512
rect 1894 2436 1994 2460
rect 527 2347 617 2393
rect 985 2347 1075 2393
rect 89 2257 135 2269
rect 89 1768 95 2257
rect 129 1768 135 2257
rect 520 2246 620 2270
rect 520 2194 544 2246
rect 596 2194 620 2246
rect 520 2170 620 2194
rect 1005 2257 1051 2269
rect 62 1744 162 1768
rect 62 1692 86 1744
rect 138 1692 162 1744
rect 62 1668 162 1692
rect 547 1681 553 2170
rect 587 1681 593 2170
rect 1005 1768 1011 2257
rect 1045 1768 1051 2257
rect 547 1669 593 1681
rect 978 1744 1078 1768
rect 978 1692 1002 1744
rect 1054 1692 1078 1744
rect 978 1668 1078 1692
rect 527 1591 617 1637
rect 985 1591 1075 1637
rect 91 1501 137 1513
rect 91 1012 97 1501
rect 131 1012 137 1501
rect 522 1490 622 1514
rect 522 1438 546 1490
rect 598 1438 622 1490
rect 522 1414 622 1438
rect 1007 1501 1053 1513
rect 64 988 164 1012
rect 64 936 88 988
rect 140 936 164 988
rect 64 912 164 936
rect 549 925 555 1414
rect 589 925 595 1414
rect 1007 1012 1013 1501
rect 1047 1012 1053 1501
rect 549 913 595 925
rect 980 988 1080 1012
rect 980 936 1004 988
rect 1056 936 1080 988
rect 980 912 1080 936
rect 527 835 617 881
rect 985 835 1075 881
rect 91 745 137 757
rect 91 256 97 745
rect 131 256 137 745
rect 522 734 622 758
rect 522 682 546 734
rect 598 682 622 734
rect 522 658 622 682
rect 1007 745 1053 757
rect 64 232 164 256
rect 64 180 88 232
rect 140 180 164 232
rect 64 156 164 180
rect 549 169 555 658
rect 589 169 595 658
rect 1007 256 1013 745
rect 1047 256 1053 745
rect 549 157 595 169
rect 980 232 1080 256
rect 980 180 1004 232
rect 1056 180 1080 232
rect 980 156 1080 180
rect 527 79 617 125
rect 985 79 1075 125
rect 1260 -40 1300 2400
rect 1443 2347 1533 2393
rect 1901 2347 1991 2393
rect 1436 2246 1536 2270
rect 1436 2194 1460 2246
rect 1512 2194 1536 2246
rect 1436 2170 1536 2194
rect 1921 2257 1967 2269
rect 1463 1681 1469 2170
rect 1503 1681 1509 2170
rect 1921 1790 1927 2257
rect 1961 1790 1967 2257
rect 2350 2246 2450 2270
rect 2350 2194 2374 2246
rect 2426 2194 2450 2246
rect 2350 2170 2450 2194
rect 2377 2160 2385 2170
rect 2417 2160 2425 2170
rect 1919 1780 1927 1790
rect 1959 1780 1967 1790
rect 1463 1669 1509 1681
rect 1892 1756 1992 1780
rect 1892 1704 1916 1756
rect 1968 1704 1992 1756
rect 1892 1680 1992 1704
rect 2379 1681 2385 2160
rect 2419 1681 2425 2160
rect 1921 1669 1967 1680
rect 2379 1669 2425 1681
rect 1443 1591 1533 1637
rect 1901 1591 1991 1637
rect 1438 1490 1538 1514
rect 1438 1438 1462 1490
rect 1514 1438 1538 1490
rect 1438 1414 1538 1438
rect 1923 1501 1969 1513
rect 1465 925 1471 1414
rect 1505 925 1511 1414
rect 1923 1034 1929 1501
rect 1963 1034 1969 1501
rect 2352 1490 2452 1514
rect 2352 1438 2376 1490
rect 2428 1438 2452 1490
rect 2352 1414 2452 1438
rect 2379 1404 2387 1414
rect 2419 1404 2427 1414
rect 1921 1024 1929 1034
rect 1961 1024 1969 1034
rect 1465 913 1511 925
rect 1894 1000 1994 1024
rect 1894 948 1918 1000
rect 1970 948 1994 1000
rect 1894 924 1994 948
rect 2381 925 2387 1404
rect 2421 925 2427 1404
rect 1923 913 1969 924
rect 2381 913 2427 925
rect 1443 835 1533 881
rect 1901 835 1991 881
rect 1438 734 1538 758
rect 1438 682 1462 734
rect 1514 682 1538 734
rect 1438 658 1538 682
rect 1923 745 1969 757
rect 1465 169 1471 658
rect 1505 169 1511 658
rect 1923 278 1929 745
rect 1963 278 1969 745
rect 2352 734 2452 758
rect 2352 682 2376 734
rect 2428 682 2452 734
rect 2352 658 2452 682
rect 2379 648 2387 658
rect 2419 648 2427 658
rect 1921 268 1929 278
rect 1961 268 1969 278
rect 1465 157 1511 169
rect 1894 244 1994 268
rect 1894 192 1918 244
rect 1970 192 1994 244
rect 1894 168 1994 192
rect 2381 169 2387 648
rect 2421 169 2427 648
rect 1923 157 1969 168
rect 2381 157 2427 169
rect 1443 79 1533 125
rect 1901 79 1991 125
<< via1 >>
rect 546 2950 598 3002
rect 1462 2950 1514 3002
rect 2376 2950 2428 3002
rect 88 2448 140 2500
rect 1004 2448 1056 2500
rect 1918 2460 1970 2512
rect 544 2194 596 2246
rect 86 1692 138 1744
rect 1002 1692 1054 1744
rect 546 1438 598 1490
rect 88 936 140 988
rect 1004 936 1056 988
rect 546 682 598 734
rect 88 180 140 232
rect 1004 180 1056 232
rect 1460 2194 1512 2246
rect 2374 2194 2426 2246
rect 1916 1704 1968 1756
rect 1462 1438 1514 1490
rect 2376 1438 2428 1490
rect 1918 948 1970 1000
rect 1462 682 1514 734
rect 2376 682 2428 734
rect 1918 192 1970 244
<< metal2 >>
rect 2352 3030 2442 3032
rect 522 3002 2442 3030
rect 522 2950 546 3002
rect 598 2950 1462 3002
rect 1514 2950 2376 3002
rect 2428 2950 2442 3002
rect 522 2916 2442 2950
rect 74 2512 1984 2546
rect 74 2500 1918 2512
rect 74 2448 88 2500
rect 140 2498 1004 2500
rect 1056 2498 1918 2500
rect 140 2448 1002 2498
rect 1058 2460 1918 2498
rect 1970 2460 1984 2512
rect 74 2442 1002 2448
rect 1058 2442 1984 2460
rect 74 2414 1984 2442
rect 1000 2410 1060 2414
rect 530 2246 2440 2292
rect 530 2194 544 2246
rect 596 2194 1460 2246
rect 1512 2194 2374 2246
rect 2426 2194 2440 2246
rect 530 2160 2440 2194
rect 72 1756 1982 1790
rect 72 1748 1916 1756
rect 72 1744 1002 1748
rect 72 1692 86 1744
rect 138 1692 1002 1744
rect 1058 1704 1916 1748
rect 1968 1704 1982 1756
rect 1058 1692 1982 1704
rect 72 1658 1982 1692
rect 532 1490 2442 1536
rect 532 1438 546 1490
rect 598 1438 1462 1490
rect 1514 1438 2376 1490
rect 2428 1438 2442 1490
rect 532 1404 2442 1438
rect 74 1000 1984 1034
rect 74 998 1918 1000
rect 74 988 1002 998
rect 74 936 88 988
rect 140 942 1002 988
rect 1058 948 1918 998
rect 1970 948 1984 1000
rect 1058 942 1984 948
rect 140 936 1004 942
rect 1056 936 1984 942
rect 74 902 1984 936
rect 532 734 2442 780
rect 532 682 546 734
rect 598 682 1462 734
rect 1514 682 2376 734
rect 2428 682 2442 734
rect 532 648 2442 682
rect 74 244 1984 278
rect 74 238 1918 244
rect 74 232 1002 238
rect 74 180 88 232
rect 140 182 1002 232
rect 1058 192 1918 238
rect 1970 192 1984 244
rect 1058 182 1984 192
rect 140 180 1004 182
rect 1056 180 1984 182
rect 74 146 1984 180
<< via2 >>
rect 1002 2448 1004 2498
rect 1004 2448 1056 2498
rect 1056 2448 1058 2498
rect 1002 2442 1058 2448
rect 1002 1744 1058 1748
rect 1002 1692 1054 1744
rect 1054 1692 1058 1744
rect 1002 988 1058 998
rect 1002 942 1004 988
rect 1004 942 1056 988
rect 1056 942 1058 988
rect 1002 232 1058 238
rect 1002 182 1004 232
rect 1004 182 1056 232
rect 1056 182 1058 232
<< metal3 >>
rect 990 2498 1070 2525
rect 990 2442 1002 2498
rect 1058 2442 1070 2498
rect 990 1748 1070 2442
rect 990 1692 1002 1748
rect 1058 1692 1070 1748
rect 990 998 1070 1692
rect 990 942 1002 998
rect 1058 942 1070 998
rect 990 238 1070 942
rect 990 182 1002 238
rect 1058 182 1070 238
rect 990 -50 1070 182
use sky130_fd_pr__nfet_01v8_lvt_USQY94  sky130_fd_pr__nfet_01v8_lvt_USQY94_0
timestamp 1663011646
transform 1 0 1259 0 1 1560
box -1302 -1603 1302 1603
<< end >>
