magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< metal4 >>
rect -651 438 651 500
rect -651 202 395 438
rect 631 202 651 438
rect -651 118 651 202
rect -651 -118 395 118
rect 631 -118 651 118
rect -651 -202 651 -118
rect -651 -438 395 -202
rect 631 -438 651 -202
rect -651 -500 651 -438
<< via4 >>
rect 395 202 631 438
rect 395 -118 631 118
rect 395 -438 631 -202
<< mimcap2 >>
rect -551 278 49 400
rect -551 -278 -369 278
rect -133 -278 49 278
rect -551 -400 49 -278
<< mimcap2contact >>
rect -369 -278 -133 278
<< metal5 >>
rect 353 438 673 501
rect -535 278 33 384
rect -535 -278 -369 278
rect -133 -278 33 278
rect -535 -384 33 -278
rect 353 202 395 438
rect 631 202 673 438
rect 353 118 673 202
rect 353 -118 395 118
rect 631 -118 673 118
rect 353 -202 673 -118
rect 353 -438 395 -202
rect 631 -438 673 -202
rect 353 -501 673 -438
<< properties >>
string FIXED_BBOX -651 -500 149 500
<< end >>
