magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -1302 -1603 1302 1603
<< nmoslvt >>
rect -1116 865 -716 1465
rect -658 865 -258 1465
rect -200 865 200 1465
rect 258 865 658 1465
rect 716 865 1116 1465
rect -1116 109 -716 709
rect -658 109 -258 709
rect -200 109 200 709
rect 258 109 658 709
rect 716 109 1116 709
rect -1116 -647 -716 -47
rect -658 -647 -258 -47
rect -200 -647 200 -47
rect 258 -647 658 -47
rect 716 -647 1116 -47
rect -1116 -1403 -716 -803
rect -658 -1403 -258 -803
rect -200 -1403 200 -803
rect 258 -1403 658 -803
rect 716 -1403 1116 -803
<< ndiff >>
rect -1174 1420 -1116 1465
rect -1174 1386 -1162 1420
rect -1128 1386 -1116 1420
rect -1174 1352 -1116 1386
rect -1174 1318 -1162 1352
rect -1128 1318 -1116 1352
rect -1174 1284 -1116 1318
rect -1174 1250 -1162 1284
rect -1128 1250 -1116 1284
rect -1174 1216 -1116 1250
rect -1174 1182 -1162 1216
rect -1128 1182 -1116 1216
rect -1174 1148 -1116 1182
rect -1174 1114 -1162 1148
rect -1128 1114 -1116 1148
rect -1174 1080 -1116 1114
rect -1174 1046 -1162 1080
rect -1128 1046 -1116 1080
rect -1174 1012 -1116 1046
rect -1174 978 -1162 1012
rect -1128 978 -1116 1012
rect -1174 944 -1116 978
rect -1174 910 -1162 944
rect -1128 910 -1116 944
rect -1174 865 -1116 910
rect -716 1420 -658 1465
rect -716 1386 -704 1420
rect -670 1386 -658 1420
rect -716 1352 -658 1386
rect -716 1318 -704 1352
rect -670 1318 -658 1352
rect -716 1284 -658 1318
rect -716 1250 -704 1284
rect -670 1250 -658 1284
rect -716 1216 -658 1250
rect -716 1182 -704 1216
rect -670 1182 -658 1216
rect -716 1148 -658 1182
rect -716 1114 -704 1148
rect -670 1114 -658 1148
rect -716 1080 -658 1114
rect -716 1046 -704 1080
rect -670 1046 -658 1080
rect -716 1012 -658 1046
rect -716 978 -704 1012
rect -670 978 -658 1012
rect -716 944 -658 978
rect -716 910 -704 944
rect -670 910 -658 944
rect -716 865 -658 910
rect -258 1420 -200 1465
rect -258 1386 -246 1420
rect -212 1386 -200 1420
rect -258 1352 -200 1386
rect -258 1318 -246 1352
rect -212 1318 -200 1352
rect -258 1284 -200 1318
rect -258 1250 -246 1284
rect -212 1250 -200 1284
rect -258 1216 -200 1250
rect -258 1182 -246 1216
rect -212 1182 -200 1216
rect -258 1148 -200 1182
rect -258 1114 -246 1148
rect -212 1114 -200 1148
rect -258 1080 -200 1114
rect -258 1046 -246 1080
rect -212 1046 -200 1080
rect -258 1012 -200 1046
rect -258 978 -246 1012
rect -212 978 -200 1012
rect -258 944 -200 978
rect -258 910 -246 944
rect -212 910 -200 944
rect -258 865 -200 910
rect 200 1420 258 1465
rect 200 1386 212 1420
rect 246 1386 258 1420
rect 200 1352 258 1386
rect 200 1318 212 1352
rect 246 1318 258 1352
rect 200 1284 258 1318
rect 200 1250 212 1284
rect 246 1250 258 1284
rect 200 1216 258 1250
rect 200 1182 212 1216
rect 246 1182 258 1216
rect 200 1148 258 1182
rect 200 1114 212 1148
rect 246 1114 258 1148
rect 200 1080 258 1114
rect 200 1046 212 1080
rect 246 1046 258 1080
rect 200 1012 258 1046
rect 200 978 212 1012
rect 246 978 258 1012
rect 200 944 258 978
rect 200 910 212 944
rect 246 910 258 944
rect 200 865 258 910
rect 658 1420 716 1465
rect 658 1386 670 1420
rect 704 1386 716 1420
rect 658 1352 716 1386
rect 658 1318 670 1352
rect 704 1318 716 1352
rect 658 1284 716 1318
rect 658 1250 670 1284
rect 704 1250 716 1284
rect 658 1216 716 1250
rect 658 1182 670 1216
rect 704 1182 716 1216
rect 658 1148 716 1182
rect 658 1114 670 1148
rect 704 1114 716 1148
rect 658 1080 716 1114
rect 658 1046 670 1080
rect 704 1046 716 1080
rect 658 1012 716 1046
rect 658 978 670 1012
rect 704 978 716 1012
rect 658 944 716 978
rect 658 910 670 944
rect 704 910 716 944
rect 658 865 716 910
rect 1116 1420 1174 1465
rect 1116 1386 1128 1420
rect 1162 1386 1174 1420
rect 1116 1352 1174 1386
rect 1116 1318 1128 1352
rect 1162 1318 1174 1352
rect 1116 1284 1174 1318
rect 1116 1250 1128 1284
rect 1162 1250 1174 1284
rect 1116 1216 1174 1250
rect 1116 1182 1128 1216
rect 1162 1182 1174 1216
rect 1116 1148 1174 1182
rect 1116 1114 1128 1148
rect 1162 1114 1174 1148
rect 1116 1080 1174 1114
rect 1116 1046 1128 1080
rect 1162 1046 1174 1080
rect 1116 1012 1174 1046
rect 1116 978 1128 1012
rect 1162 978 1174 1012
rect 1116 944 1174 978
rect 1116 910 1128 944
rect 1162 910 1174 944
rect 1116 865 1174 910
rect -1174 664 -1116 709
rect -1174 630 -1162 664
rect -1128 630 -1116 664
rect -1174 596 -1116 630
rect -1174 562 -1162 596
rect -1128 562 -1116 596
rect -1174 528 -1116 562
rect -1174 494 -1162 528
rect -1128 494 -1116 528
rect -1174 460 -1116 494
rect -1174 426 -1162 460
rect -1128 426 -1116 460
rect -1174 392 -1116 426
rect -1174 358 -1162 392
rect -1128 358 -1116 392
rect -1174 324 -1116 358
rect -1174 290 -1162 324
rect -1128 290 -1116 324
rect -1174 256 -1116 290
rect -1174 222 -1162 256
rect -1128 222 -1116 256
rect -1174 188 -1116 222
rect -1174 154 -1162 188
rect -1128 154 -1116 188
rect -1174 109 -1116 154
rect -716 664 -658 709
rect -716 630 -704 664
rect -670 630 -658 664
rect -716 596 -658 630
rect -716 562 -704 596
rect -670 562 -658 596
rect -716 528 -658 562
rect -716 494 -704 528
rect -670 494 -658 528
rect -716 460 -658 494
rect -716 426 -704 460
rect -670 426 -658 460
rect -716 392 -658 426
rect -716 358 -704 392
rect -670 358 -658 392
rect -716 324 -658 358
rect -716 290 -704 324
rect -670 290 -658 324
rect -716 256 -658 290
rect -716 222 -704 256
rect -670 222 -658 256
rect -716 188 -658 222
rect -716 154 -704 188
rect -670 154 -658 188
rect -716 109 -658 154
rect -258 664 -200 709
rect -258 630 -246 664
rect -212 630 -200 664
rect -258 596 -200 630
rect -258 562 -246 596
rect -212 562 -200 596
rect -258 528 -200 562
rect -258 494 -246 528
rect -212 494 -200 528
rect -258 460 -200 494
rect -258 426 -246 460
rect -212 426 -200 460
rect -258 392 -200 426
rect -258 358 -246 392
rect -212 358 -200 392
rect -258 324 -200 358
rect -258 290 -246 324
rect -212 290 -200 324
rect -258 256 -200 290
rect -258 222 -246 256
rect -212 222 -200 256
rect -258 188 -200 222
rect -258 154 -246 188
rect -212 154 -200 188
rect -258 109 -200 154
rect 200 664 258 709
rect 200 630 212 664
rect 246 630 258 664
rect 200 596 258 630
rect 200 562 212 596
rect 246 562 258 596
rect 200 528 258 562
rect 200 494 212 528
rect 246 494 258 528
rect 200 460 258 494
rect 200 426 212 460
rect 246 426 258 460
rect 200 392 258 426
rect 200 358 212 392
rect 246 358 258 392
rect 200 324 258 358
rect 200 290 212 324
rect 246 290 258 324
rect 200 256 258 290
rect 200 222 212 256
rect 246 222 258 256
rect 200 188 258 222
rect 200 154 212 188
rect 246 154 258 188
rect 200 109 258 154
rect 658 664 716 709
rect 658 630 670 664
rect 704 630 716 664
rect 658 596 716 630
rect 658 562 670 596
rect 704 562 716 596
rect 658 528 716 562
rect 658 494 670 528
rect 704 494 716 528
rect 658 460 716 494
rect 658 426 670 460
rect 704 426 716 460
rect 658 392 716 426
rect 658 358 670 392
rect 704 358 716 392
rect 658 324 716 358
rect 658 290 670 324
rect 704 290 716 324
rect 658 256 716 290
rect 658 222 670 256
rect 704 222 716 256
rect 658 188 716 222
rect 658 154 670 188
rect 704 154 716 188
rect 658 109 716 154
rect 1116 664 1174 709
rect 1116 630 1128 664
rect 1162 630 1174 664
rect 1116 596 1174 630
rect 1116 562 1128 596
rect 1162 562 1174 596
rect 1116 528 1174 562
rect 1116 494 1128 528
rect 1162 494 1174 528
rect 1116 460 1174 494
rect 1116 426 1128 460
rect 1162 426 1174 460
rect 1116 392 1174 426
rect 1116 358 1128 392
rect 1162 358 1174 392
rect 1116 324 1174 358
rect 1116 290 1128 324
rect 1162 290 1174 324
rect 1116 256 1174 290
rect 1116 222 1128 256
rect 1162 222 1174 256
rect 1116 188 1174 222
rect 1116 154 1128 188
rect 1162 154 1174 188
rect 1116 109 1174 154
rect -1174 -92 -1116 -47
rect -1174 -126 -1162 -92
rect -1128 -126 -1116 -92
rect -1174 -160 -1116 -126
rect -1174 -194 -1162 -160
rect -1128 -194 -1116 -160
rect -1174 -228 -1116 -194
rect -1174 -262 -1162 -228
rect -1128 -262 -1116 -228
rect -1174 -296 -1116 -262
rect -1174 -330 -1162 -296
rect -1128 -330 -1116 -296
rect -1174 -364 -1116 -330
rect -1174 -398 -1162 -364
rect -1128 -398 -1116 -364
rect -1174 -432 -1116 -398
rect -1174 -466 -1162 -432
rect -1128 -466 -1116 -432
rect -1174 -500 -1116 -466
rect -1174 -534 -1162 -500
rect -1128 -534 -1116 -500
rect -1174 -568 -1116 -534
rect -1174 -602 -1162 -568
rect -1128 -602 -1116 -568
rect -1174 -647 -1116 -602
rect -716 -92 -658 -47
rect -716 -126 -704 -92
rect -670 -126 -658 -92
rect -716 -160 -658 -126
rect -716 -194 -704 -160
rect -670 -194 -658 -160
rect -716 -228 -658 -194
rect -716 -262 -704 -228
rect -670 -262 -658 -228
rect -716 -296 -658 -262
rect -716 -330 -704 -296
rect -670 -330 -658 -296
rect -716 -364 -658 -330
rect -716 -398 -704 -364
rect -670 -398 -658 -364
rect -716 -432 -658 -398
rect -716 -466 -704 -432
rect -670 -466 -658 -432
rect -716 -500 -658 -466
rect -716 -534 -704 -500
rect -670 -534 -658 -500
rect -716 -568 -658 -534
rect -716 -602 -704 -568
rect -670 -602 -658 -568
rect -716 -647 -658 -602
rect -258 -92 -200 -47
rect -258 -126 -246 -92
rect -212 -126 -200 -92
rect -258 -160 -200 -126
rect -258 -194 -246 -160
rect -212 -194 -200 -160
rect -258 -228 -200 -194
rect -258 -262 -246 -228
rect -212 -262 -200 -228
rect -258 -296 -200 -262
rect -258 -330 -246 -296
rect -212 -330 -200 -296
rect -258 -364 -200 -330
rect -258 -398 -246 -364
rect -212 -398 -200 -364
rect -258 -432 -200 -398
rect -258 -466 -246 -432
rect -212 -466 -200 -432
rect -258 -500 -200 -466
rect -258 -534 -246 -500
rect -212 -534 -200 -500
rect -258 -568 -200 -534
rect -258 -602 -246 -568
rect -212 -602 -200 -568
rect -258 -647 -200 -602
rect 200 -92 258 -47
rect 200 -126 212 -92
rect 246 -126 258 -92
rect 200 -160 258 -126
rect 200 -194 212 -160
rect 246 -194 258 -160
rect 200 -228 258 -194
rect 200 -262 212 -228
rect 246 -262 258 -228
rect 200 -296 258 -262
rect 200 -330 212 -296
rect 246 -330 258 -296
rect 200 -364 258 -330
rect 200 -398 212 -364
rect 246 -398 258 -364
rect 200 -432 258 -398
rect 200 -466 212 -432
rect 246 -466 258 -432
rect 200 -500 258 -466
rect 200 -534 212 -500
rect 246 -534 258 -500
rect 200 -568 258 -534
rect 200 -602 212 -568
rect 246 -602 258 -568
rect 200 -647 258 -602
rect 658 -92 716 -47
rect 658 -126 670 -92
rect 704 -126 716 -92
rect 658 -160 716 -126
rect 658 -194 670 -160
rect 704 -194 716 -160
rect 658 -228 716 -194
rect 658 -262 670 -228
rect 704 -262 716 -228
rect 658 -296 716 -262
rect 658 -330 670 -296
rect 704 -330 716 -296
rect 658 -364 716 -330
rect 658 -398 670 -364
rect 704 -398 716 -364
rect 658 -432 716 -398
rect 658 -466 670 -432
rect 704 -466 716 -432
rect 658 -500 716 -466
rect 658 -534 670 -500
rect 704 -534 716 -500
rect 658 -568 716 -534
rect 658 -602 670 -568
rect 704 -602 716 -568
rect 658 -647 716 -602
rect 1116 -92 1174 -47
rect 1116 -126 1128 -92
rect 1162 -126 1174 -92
rect 1116 -160 1174 -126
rect 1116 -194 1128 -160
rect 1162 -194 1174 -160
rect 1116 -228 1174 -194
rect 1116 -262 1128 -228
rect 1162 -262 1174 -228
rect 1116 -296 1174 -262
rect 1116 -330 1128 -296
rect 1162 -330 1174 -296
rect 1116 -364 1174 -330
rect 1116 -398 1128 -364
rect 1162 -398 1174 -364
rect 1116 -432 1174 -398
rect 1116 -466 1128 -432
rect 1162 -466 1174 -432
rect 1116 -500 1174 -466
rect 1116 -534 1128 -500
rect 1162 -534 1174 -500
rect 1116 -568 1174 -534
rect 1116 -602 1128 -568
rect 1162 -602 1174 -568
rect 1116 -647 1174 -602
rect -1174 -848 -1116 -803
rect -1174 -882 -1162 -848
rect -1128 -882 -1116 -848
rect -1174 -916 -1116 -882
rect -1174 -950 -1162 -916
rect -1128 -950 -1116 -916
rect -1174 -984 -1116 -950
rect -1174 -1018 -1162 -984
rect -1128 -1018 -1116 -984
rect -1174 -1052 -1116 -1018
rect -1174 -1086 -1162 -1052
rect -1128 -1086 -1116 -1052
rect -1174 -1120 -1116 -1086
rect -1174 -1154 -1162 -1120
rect -1128 -1154 -1116 -1120
rect -1174 -1188 -1116 -1154
rect -1174 -1222 -1162 -1188
rect -1128 -1222 -1116 -1188
rect -1174 -1256 -1116 -1222
rect -1174 -1290 -1162 -1256
rect -1128 -1290 -1116 -1256
rect -1174 -1324 -1116 -1290
rect -1174 -1358 -1162 -1324
rect -1128 -1358 -1116 -1324
rect -1174 -1403 -1116 -1358
rect -716 -848 -658 -803
rect -716 -882 -704 -848
rect -670 -882 -658 -848
rect -716 -916 -658 -882
rect -716 -950 -704 -916
rect -670 -950 -658 -916
rect -716 -984 -658 -950
rect -716 -1018 -704 -984
rect -670 -1018 -658 -984
rect -716 -1052 -658 -1018
rect -716 -1086 -704 -1052
rect -670 -1086 -658 -1052
rect -716 -1120 -658 -1086
rect -716 -1154 -704 -1120
rect -670 -1154 -658 -1120
rect -716 -1188 -658 -1154
rect -716 -1222 -704 -1188
rect -670 -1222 -658 -1188
rect -716 -1256 -658 -1222
rect -716 -1290 -704 -1256
rect -670 -1290 -658 -1256
rect -716 -1324 -658 -1290
rect -716 -1358 -704 -1324
rect -670 -1358 -658 -1324
rect -716 -1403 -658 -1358
rect -258 -848 -200 -803
rect -258 -882 -246 -848
rect -212 -882 -200 -848
rect -258 -916 -200 -882
rect -258 -950 -246 -916
rect -212 -950 -200 -916
rect -258 -984 -200 -950
rect -258 -1018 -246 -984
rect -212 -1018 -200 -984
rect -258 -1052 -200 -1018
rect -258 -1086 -246 -1052
rect -212 -1086 -200 -1052
rect -258 -1120 -200 -1086
rect -258 -1154 -246 -1120
rect -212 -1154 -200 -1120
rect -258 -1188 -200 -1154
rect -258 -1222 -246 -1188
rect -212 -1222 -200 -1188
rect -258 -1256 -200 -1222
rect -258 -1290 -246 -1256
rect -212 -1290 -200 -1256
rect -258 -1324 -200 -1290
rect -258 -1358 -246 -1324
rect -212 -1358 -200 -1324
rect -258 -1403 -200 -1358
rect 200 -848 258 -803
rect 200 -882 212 -848
rect 246 -882 258 -848
rect 200 -916 258 -882
rect 200 -950 212 -916
rect 246 -950 258 -916
rect 200 -984 258 -950
rect 200 -1018 212 -984
rect 246 -1018 258 -984
rect 200 -1052 258 -1018
rect 200 -1086 212 -1052
rect 246 -1086 258 -1052
rect 200 -1120 258 -1086
rect 200 -1154 212 -1120
rect 246 -1154 258 -1120
rect 200 -1188 258 -1154
rect 200 -1222 212 -1188
rect 246 -1222 258 -1188
rect 200 -1256 258 -1222
rect 200 -1290 212 -1256
rect 246 -1290 258 -1256
rect 200 -1324 258 -1290
rect 200 -1358 212 -1324
rect 246 -1358 258 -1324
rect 200 -1403 258 -1358
rect 658 -848 716 -803
rect 658 -882 670 -848
rect 704 -882 716 -848
rect 658 -916 716 -882
rect 658 -950 670 -916
rect 704 -950 716 -916
rect 658 -984 716 -950
rect 658 -1018 670 -984
rect 704 -1018 716 -984
rect 658 -1052 716 -1018
rect 658 -1086 670 -1052
rect 704 -1086 716 -1052
rect 658 -1120 716 -1086
rect 658 -1154 670 -1120
rect 704 -1154 716 -1120
rect 658 -1188 716 -1154
rect 658 -1222 670 -1188
rect 704 -1222 716 -1188
rect 658 -1256 716 -1222
rect 658 -1290 670 -1256
rect 704 -1290 716 -1256
rect 658 -1324 716 -1290
rect 658 -1358 670 -1324
rect 704 -1358 716 -1324
rect 658 -1403 716 -1358
rect 1116 -848 1174 -803
rect 1116 -882 1128 -848
rect 1162 -882 1174 -848
rect 1116 -916 1174 -882
rect 1116 -950 1128 -916
rect 1162 -950 1174 -916
rect 1116 -984 1174 -950
rect 1116 -1018 1128 -984
rect 1162 -1018 1174 -984
rect 1116 -1052 1174 -1018
rect 1116 -1086 1128 -1052
rect 1162 -1086 1174 -1052
rect 1116 -1120 1174 -1086
rect 1116 -1154 1128 -1120
rect 1162 -1154 1174 -1120
rect 1116 -1188 1174 -1154
rect 1116 -1222 1128 -1188
rect 1162 -1222 1174 -1188
rect 1116 -1256 1174 -1222
rect 1116 -1290 1128 -1256
rect 1162 -1290 1174 -1256
rect 1116 -1324 1174 -1290
rect 1116 -1358 1128 -1324
rect 1162 -1358 1174 -1324
rect 1116 -1403 1174 -1358
<< ndiffc >>
rect -1162 1386 -1128 1420
rect -1162 1318 -1128 1352
rect -1162 1250 -1128 1284
rect -1162 1182 -1128 1216
rect -1162 1114 -1128 1148
rect -1162 1046 -1128 1080
rect -1162 978 -1128 1012
rect -1162 910 -1128 944
rect -704 1386 -670 1420
rect -704 1318 -670 1352
rect -704 1250 -670 1284
rect -704 1182 -670 1216
rect -704 1114 -670 1148
rect -704 1046 -670 1080
rect -704 978 -670 1012
rect -704 910 -670 944
rect -246 1386 -212 1420
rect -246 1318 -212 1352
rect -246 1250 -212 1284
rect -246 1182 -212 1216
rect -246 1114 -212 1148
rect -246 1046 -212 1080
rect -246 978 -212 1012
rect -246 910 -212 944
rect 212 1386 246 1420
rect 212 1318 246 1352
rect 212 1250 246 1284
rect 212 1182 246 1216
rect 212 1114 246 1148
rect 212 1046 246 1080
rect 212 978 246 1012
rect 212 910 246 944
rect 670 1386 704 1420
rect 670 1318 704 1352
rect 670 1250 704 1284
rect 670 1182 704 1216
rect 670 1114 704 1148
rect 670 1046 704 1080
rect 670 978 704 1012
rect 670 910 704 944
rect 1128 1386 1162 1420
rect 1128 1318 1162 1352
rect 1128 1250 1162 1284
rect 1128 1182 1162 1216
rect 1128 1114 1162 1148
rect 1128 1046 1162 1080
rect 1128 978 1162 1012
rect 1128 910 1162 944
rect -1162 630 -1128 664
rect -1162 562 -1128 596
rect -1162 494 -1128 528
rect -1162 426 -1128 460
rect -1162 358 -1128 392
rect -1162 290 -1128 324
rect -1162 222 -1128 256
rect -1162 154 -1128 188
rect -704 630 -670 664
rect -704 562 -670 596
rect -704 494 -670 528
rect -704 426 -670 460
rect -704 358 -670 392
rect -704 290 -670 324
rect -704 222 -670 256
rect -704 154 -670 188
rect -246 630 -212 664
rect -246 562 -212 596
rect -246 494 -212 528
rect -246 426 -212 460
rect -246 358 -212 392
rect -246 290 -212 324
rect -246 222 -212 256
rect -246 154 -212 188
rect 212 630 246 664
rect 212 562 246 596
rect 212 494 246 528
rect 212 426 246 460
rect 212 358 246 392
rect 212 290 246 324
rect 212 222 246 256
rect 212 154 246 188
rect 670 630 704 664
rect 670 562 704 596
rect 670 494 704 528
rect 670 426 704 460
rect 670 358 704 392
rect 670 290 704 324
rect 670 222 704 256
rect 670 154 704 188
rect 1128 630 1162 664
rect 1128 562 1162 596
rect 1128 494 1162 528
rect 1128 426 1162 460
rect 1128 358 1162 392
rect 1128 290 1162 324
rect 1128 222 1162 256
rect 1128 154 1162 188
rect -1162 -126 -1128 -92
rect -1162 -194 -1128 -160
rect -1162 -262 -1128 -228
rect -1162 -330 -1128 -296
rect -1162 -398 -1128 -364
rect -1162 -466 -1128 -432
rect -1162 -534 -1128 -500
rect -1162 -602 -1128 -568
rect -704 -126 -670 -92
rect -704 -194 -670 -160
rect -704 -262 -670 -228
rect -704 -330 -670 -296
rect -704 -398 -670 -364
rect -704 -466 -670 -432
rect -704 -534 -670 -500
rect -704 -602 -670 -568
rect -246 -126 -212 -92
rect -246 -194 -212 -160
rect -246 -262 -212 -228
rect -246 -330 -212 -296
rect -246 -398 -212 -364
rect -246 -466 -212 -432
rect -246 -534 -212 -500
rect -246 -602 -212 -568
rect 212 -126 246 -92
rect 212 -194 246 -160
rect 212 -262 246 -228
rect 212 -330 246 -296
rect 212 -398 246 -364
rect 212 -466 246 -432
rect 212 -534 246 -500
rect 212 -602 246 -568
rect 670 -126 704 -92
rect 670 -194 704 -160
rect 670 -262 704 -228
rect 670 -330 704 -296
rect 670 -398 704 -364
rect 670 -466 704 -432
rect 670 -534 704 -500
rect 670 -602 704 -568
rect 1128 -126 1162 -92
rect 1128 -194 1162 -160
rect 1128 -262 1162 -228
rect 1128 -330 1162 -296
rect 1128 -398 1162 -364
rect 1128 -466 1162 -432
rect 1128 -534 1162 -500
rect 1128 -602 1162 -568
rect -1162 -882 -1128 -848
rect -1162 -950 -1128 -916
rect -1162 -1018 -1128 -984
rect -1162 -1086 -1128 -1052
rect -1162 -1154 -1128 -1120
rect -1162 -1222 -1128 -1188
rect -1162 -1290 -1128 -1256
rect -1162 -1358 -1128 -1324
rect -704 -882 -670 -848
rect -704 -950 -670 -916
rect -704 -1018 -670 -984
rect -704 -1086 -670 -1052
rect -704 -1154 -670 -1120
rect -704 -1222 -670 -1188
rect -704 -1290 -670 -1256
rect -704 -1358 -670 -1324
rect -246 -882 -212 -848
rect -246 -950 -212 -916
rect -246 -1018 -212 -984
rect -246 -1086 -212 -1052
rect -246 -1154 -212 -1120
rect -246 -1222 -212 -1188
rect -246 -1290 -212 -1256
rect -246 -1358 -212 -1324
rect 212 -882 246 -848
rect 212 -950 246 -916
rect 212 -1018 246 -984
rect 212 -1086 246 -1052
rect 212 -1154 246 -1120
rect 212 -1222 246 -1188
rect 212 -1290 246 -1256
rect 212 -1358 246 -1324
rect 670 -882 704 -848
rect 670 -950 704 -916
rect 670 -1018 704 -984
rect 670 -1086 704 -1052
rect 670 -1154 704 -1120
rect 670 -1222 704 -1188
rect 670 -1290 704 -1256
rect 670 -1358 704 -1324
rect 1128 -882 1162 -848
rect 1128 -950 1162 -916
rect 1128 -1018 1162 -984
rect 1128 -1086 1162 -1052
rect 1128 -1154 1162 -1120
rect 1128 -1222 1162 -1188
rect 1128 -1290 1162 -1256
rect 1128 -1358 1162 -1324
<< psubdiff >>
rect -1276 1543 -1173 1577
rect -1139 1543 -1105 1577
rect -1071 1543 -1037 1577
rect -1003 1543 -969 1577
rect -935 1543 -901 1577
rect -867 1543 -833 1577
rect -799 1543 -765 1577
rect -731 1543 -697 1577
rect -663 1543 -629 1577
rect -595 1543 -561 1577
rect -527 1543 -493 1577
rect -459 1543 -425 1577
rect -391 1543 -357 1577
rect -323 1543 -289 1577
rect -255 1543 -221 1577
rect -187 1543 -153 1577
rect -119 1543 -85 1577
rect -51 1543 -17 1577
rect 17 1543 51 1577
rect 85 1543 119 1577
rect 153 1543 187 1577
rect 221 1543 255 1577
rect 289 1543 323 1577
rect 357 1543 391 1577
rect 425 1543 459 1577
rect 493 1543 527 1577
rect 561 1543 595 1577
rect 629 1543 663 1577
rect 697 1543 731 1577
rect 765 1543 799 1577
rect 833 1543 867 1577
rect 901 1543 935 1577
rect 969 1543 1003 1577
rect 1037 1543 1071 1577
rect 1105 1543 1139 1577
rect 1173 1543 1276 1577
rect -1276 -1543 -1242 1543
rect 1242 -1543 1276 1543
rect -1276 -1577 -1173 -1543
rect -1139 -1577 -1105 -1543
rect -1071 -1577 -1037 -1543
rect -1003 -1577 -969 -1543
rect -935 -1577 -901 -1543
rect -867 -1577 -833 -1543
rect -799 -1577 -765 -1543
rect -731 -1577 -697 -1543
rect -663 -1577 -629 -1543
rect -595 -1577 -561 -1543
rect -527 -1577 -493 -1543
rect -459 -1577 -425 -1543
rect -391 -1577 -357 -1543
rect -323 -1577 -289 -1543
rect -255 -1577 -221 -1543
rect -187 -1577 -153 -1543
rect -119 -1577 -85 -1543
rect -51 -1577 -17 -1543
rect 17 -1577 51 -1543
rect 85 -1577 119 -1543
rect 153 -1577 187 -1543
rect 221 -1577 255 -1543
rect 289 -1577 323 -1543
rect 357 -1577 391 -1543
rect 425 -1577 459 -1543
rect 493 -1577 527 -1543
rect 561 -1577 595 -1543
rect 629 -1577 663 -1543
rect 697 -1577 731 -1543
rect 765 -1577 799 -1543
rect 833 -1577 867 -1543
rect 901 -1577 935 -1543
rect 969 -1577 1003 -1543
rect 1037 -1577 1071 -1543
rect 1105 -1577 1139 -1543
rect 1173 -1577 1276 -1543
<< psubdiffcont >>
rect -1173 1543 -1139 1577
rect -1105 1543 -1071 1577
rect -1037 1543 -1003 1577
rect -969 1543 -935 1577
rect -901 1543 -867 1577
rect -833 1543 -799 1577
rect -765 1543 -731 1577
rect -697 1543 -663 1577
rect -629 1543 -595 1577
rect -561 1543 -527 1577
rect -493 1543 -459 1577
rect -425 1543 -391 1577
rect -357 1543 -323 1577
rect -289 1543 -255 1577
rect -221 1543 -187 1577
rect -153 1543 -119 1577
rect -85 1543 -51 1577
rect -17 1543 17 1577
rect 51 1543 85 1577
rect 119 1543 153 1577
rect 187 1543 221 1577
rect 255 1543 289 1577
rect 323 1543 357 1577
rect 391 1543 425 1577
rect 459 1543 493 1577
rect 527 1543 561 1577
rect 595 1543 629 1577
rect 663 1543 697 1577
rect 731 1543 765 1577
rect 799 1543 833 1577
rect 867 1543 901 1577
rect 935 1543 969 1577
rect 1003 1543 1037 1577
rect 1071 1543 1105 1577
rect 1139 1543 1173 1577
rect -1173 -1577 -1139 -1543
rect -1105 -1577 -1071 -1543
rect -1037 -1577 -1003 -1543
rect -969 -1577 -935 -1543
rect -901 -1577 -867 -1543
rect -833 -1577 -799 -1543
rect -765 -1577 -731 -1543
rect -697 -1577 -663 -1543
rect -629 -1577 -595 -1543
rect -561 -1577 -527 -1543
rect -493 -1577 -459 -1543
rect -425 -1577 -391 -1543
rect -357 -1577 -323 -1543
rect -289 -1577 -255 -1543
rect -221 -1577 -187 -1543
rect -153 -1577 -119 -1543
rect -85 -1577 -51 -1543
rect -17 -1577 17 -1543
rect 51 -1577 85 -1543
rect 119 -1577 153 -1543
rect 187 -1577 221 -1543
rect 255 -1577 289 -1543
rect 323 -1577 357 -1543
rect 391 -1577 425 -1543
rect 459 -1577 493 -1543
rect 527 -1577 561 -1543
rect 595 -1577 629 -1543
rect 663 -1577 697 -1543
rect 731 -1577 765 -1543
rect 799 -1577 833 -1543
rect 867 -1577 901 -1543
rect 935 -1577 969 -1543
rect 1003 -1577 1037 -1543
rect 1071 -1577 1105 -1543
rect 1139 -1577 1173 -1543
<< poly >>
rect -1116 1465 -716 1491
rect -658 1465 -258 1491
rect -200 1465 200 1491
rect 258 1465 658 1491
rect 716 1465 1116 1491
rect -1116 827 -716 865
rect -1116 793 -1069 827
rect -1035 793 -1001 827
rect -967 793 -933 827
rect -899 793 -865 827
rect -831 793 -797 827
rect -763 793 -716 827
rect -1116 777 -716 793
rect -658 827 -258 865
rect -658 793 -611 827
rect -577 793 -543 827
rect -509 793 -475 827
rect -441 793 -407 827
rect -373 793 -339 827
rect -305 793 -258 827
rect -658 777 -258 793
rect -200 827 200 865
rect -200 793 -153 827
rect -119 793 -85 827
rect -51 793 -17 827
rect 17 793 51 827
rect 85 793 119 827
rect 153 793 200 827
rect -200 777 200 793
rect 258 827 658 865
rect 258 793 305 827
rect 339 793 373 827
rect 407 793 441 827
rect 475 793 509 827
rect 543 793 577 827
rect 611 793 658 827
rect 258 777 658 793
rect 716 827 1116 865
rect 716 793 763 827
rect 797 793 831 827
rect 865 793 899 827
rect 933 793 967 827
rect 1001 793 1035 827
rect 1069 793 1116 827
rect 716 777 1116 793
rect -1116 709 -716 735
rect -658 709 -258 735
rect -200 709 200 735
rect 258 709 658 735
rect 716 709 1116 735
rect -1116 71 -716 109
rect -1116 37 -1069 71
rect -1035 37 -1001 71
rect -967 37 -933 71
rect -899 37 -865 71
rect -831 37 -797 71
rect -763 37 -716 71
rect -1116 21 -716 37
rect -658 71 -258 109
rect -658 37 -611 71
rect -577 37 -543 71
rect -509 37 -475 71
rect -441 37 -407 71
rect -373 37 -339 71
rect -305 37 -258 71
rect -658 21 -258 37
rect -200 71 200 109
rect -200 37 -153 71
rect -119 37 -85 71
rect -51 37 -17 71
rect 17 37 51 71
rect 85 37 119 71
rect 153 37 200 71
rect -200 21 200 37
rect 258 71 658 109
rect 258 37 305 71
rect 339 37 373 71
rect 407 37 441 71
rect 475 37 509 71
rect 543 37 577 71
rect 611 37 658 71
rect 258 21 658 37
rect 716 71 1116 109
rect 716 37 763 71
rect 797 37 831 71
rect 865 37 899 71
rect 933 37 967 71
rect 1001 37 1035 71
rect 1069 37 1116 71
rect 716 21 1116 37
rect -1116 -47 -716 -21
rect -658 -47 -258 -21
rect -200 -47 200 -21
rect 258 -47 658 -21
rect 716 -47 1116 -21
rect -1116 -685 -716 -647
rect -1116 -719 -1069 -685
rect -1035 -719 -1001 -685
rect -967 -719 -933 -685
rect -899 -719 -865 -685
rect -831 -719 -797 -685
rect -763 -719 -716 -685
rect -1116 -735 -716 -719
rect -658 -685 -258 -647
rect -658 -719 -611 -685
rect -577 -719 -543 -685
rect -509 -719 -475 -685
rect -441 -719 -407 -685
rect -373 -719 -339 -685
rect -305 -719 -258 -685
rect -658 -735 -258 -719
rect -200 -685 200 -647
rect -200 -719 -153 -685
rect -119 -719 -85 -685
rect -51 -719 -17 -685
rect 17 -719 51 -685
rect 85 -719 119 -685
rect 153 -719 200 -685
rect -200 -735 200 -719
rect 258 -685 658 -647
rect 258 -719 305 -685
rect 339 -719 373 -685
rect 407 -719 441 -685
rect 475 -719 509 -685
rect 543 -719 577 -685
rect 611 -719 658 -685
rect 258 -735 658 -719
rect 716 -685 1116 -647
rect 716 -719 763 -685
rect 797 -719 831 -685
rect 865 -719 899 -685
rect 933 -719 967 -685
rect 1001 -719 1035 -685
rect 1069 -719 1116 -685
rect 716 -735 1116 -719
rect -1116 -803 -716 -777
rect -658 -803 -258 -777
rect -200 -803 200 -777
rect 258 -803 658 -777
rect 716 -803 1116 -777
rect -1116 -1441 -716 -1403
rect -1116 -1475 -1069 -1441
rect -1035 -1475 -1001 -1441
rect -967 -1475 -933 -1441
rect -899 -1475 -865 -1441
rect -831 -1475 -797 -1441
rect -763 -1475 -716 -1441
rect -1116 -1491 -716 -1475
rect -658 -1441 -258 -1403
rect -658 -1475 -611 -1441
rect -577 -1475 -543 -1441
rect -509 -1475 -475 -1441
rect -441 -1475 -407 -1441
rect -373 -1475 -339 -1441
rect -305 -1475 -258 -1441
rect -658 -1491 -258 -1475
rect -200 -1441 200 -1403
rect -200 -1475 -153 -1441
rect -119 -1475 -85 -1441
rect -51 -1475 -17 -1441
rect 17 -1475 51 -1441
rect 85 -1475 119 -1441
rect 153 -1475 200 -1441
rect -200 -1491 200 -1475
rect 258 -1441 658 -1403
rect 258 -1475 305 -1441
rect 339 -1475 373 -1441
rect 407 -1475 441 -1441
rect 475 -1475 509 -1441
rect 543 -1475 577 -1441
rect 611 -1475 658 -1441
rect 258 -1491 658 -1475
rect 716 -1441 1116 -1403
rect 716 -1475 763 -1441
rect 797 -1475 831 -1441
rect 865 -1475 899 -1441
rect 933 -1475 967 -1441
rect 1001 -1475 1035 -1441
rect 1069 -1475 1116 -1441
rect 716 -1491 1116 -1475
<< polycont >>
rect -1069 793 -1035 827
rect -1001 793 -967 827
rect -933 793 -899 827
rect -865 793 -831 827
rect -797 793 -763 827
rect -611 793 -577 827
rect -543 793 -509 827
rect -475 793 -441 827
rect -407 793 -373 827
rect -339 793 -305 827
rect -153 793 -119 827
rect -85 793 -51 827
rect -17 793 17 827
rect 51 793 85 827
rect 119 793 153 827
rect 305 793 339 827
rect 373 793 407 827
rect 441 793 475 827
rect 509 793 543 827
rect 577 793 611 827
rect 763 793 797 827
rect 831 793 865 827
rect 899 793 933 827
rect 967 793 1001 827
rect 1035 793 1069 827
rect -1069 37 -1035 71
rect -1001 37 -967 71
rect -933 37 -899 71
rect -865 37 -831 71
rect -797 37 -763 71
rect -611 37 -577 71
rect -543 37 -509 71
rect -475 37 -441 71
rect -407 37 -373 71
rect -339 37 -305 71
rect -153 37 -119 71
rect -85 37 -51 71
rect -17 37 17 71
rect 51 37 85 71
rect 119 37 153 71
rect 305 37 339 71
rect 373 37 407 71
rect 441 37 475 71
rect 509 37 543 71
rect 577 37 611 71
rect 763 37 797 71
rect 831 37 865 71
rect 899 37 933 71
rect 967 37 1001 71
rect 1035 37 1069 71
rect -1069 -719 -1035 -685
rect -1001 -719 -967 -685
rect -933 -719 -899 -685
rect -865 -719 -831 -685
rect -797 -719 -763 -685
rect -611 -719 -577 -685
rect -543 -719 -509 -685
rect -475 -719 -441 -685
rect -407 -719 -373 -685
rect -339 -719 -305 -685
rect -153 -719 -119 -685
rect -85 -719 -51 -685
rect -17 -719 17 -685
rect 51 -719 85 -685
rect 119 -719 153 -685
rect 305 -719 339 -685
rect 373 -719 407 -685
rect 441 -719 475 -685
rect 509 -719 543 -685
rect 577 -719 611 -685
rect 763 -719 797 -685
rect 831 -719 865 -685
rect 899 -719 933 -685
rect 967 -719 1001 -685
rect 1035 -719 1069 -685
rect -1069 -1475 -1035 -1441
rect -1001 -1475 -967 -1441
rect -933 -1475 -899 -1441
rect -865 -1475 -831 -1441
rect -797 -1475 -763 -1441
rect -611 -1475 -577 -1441
rect -543 -1475 -509 -1441
rect -475 -1475 -441 -1441
rect -407 -1475 -373 -1441
rect -339 -1475 -305 -1441
rect -153 -1475 -119 -1441
rect -85 -1475 -51 -1441
rect -17 -1475 17 -1441
rect 51 -1475 85 -1441
rect 119 -1475 153 -1441
rect 305 -1475 339 -1441
rect 373 -1475 407 -1441
rect 441 -1475 475 -1441
rect 509 -1475 543 -1441
rect 577 -1475 611 -1441
rect 763 -1475 797 -1441
rect 831 -1475 865 -1441
rect 899 -1475 933 -1441
rect 967 -1475 1001 -1441
rect 1035 -1475 1069 -1441
<< locali >>
rect -1276 1543 -1173 1577
rect -1139 1543 -1105 1577
rect -1071 1543 -1037 1577
rect -1003 1543 -969 1577
rect -935 1543 -901 1577
rect -867 1543 -833 1577
rect -799 1543 -765 1577
rect -731 1543 -697 1577
rect -663 1543 -629 1577
rect -595 1543 -561 1577
rect -527 1543 -493 1577
rect -459 1543 -425 1577
rect -391 1543 -357 1577
rect -323 1543 -289 1577
rect -255 1543 -221 1577
rect -187 1543 -153 1577
rect -119 1543 -85 1577
rect -51 1543 -17 1577
rect 17 1543 51 1577
rect 85 1543 119 1577
rect 153 1543 187 1577
rect 221 1543 255 1577
rect 289 1543 323 1577
rect 357 1543 391 1577
rect 425 1543 459 1577
rect 493 1543 527 1577
rect 561 1543 595 1577
rect 629 1543 663 1577
rect 697 1543 731 1577
rect 765 1543 799 1577
rect 833 1543 867 1577
rect 901 1543 935 1577
rect 969 1543 1003 1577
rect 1037 1543 1071 1577
rect 1105 1543 1139 1577
rect 1173 1543 1276 1577
rect -1276 -1543 -1242 1543
rect -1162 1434 -1128 1469
rect -1162 1362 -1128 1386
rect -1162 1290 -1128 1318
rect -1162 1218 -1128 1250
rect -1162 1148 -1128 1182
rect -1162 1080 -1128 1112
rect -1162 1012 -1128 1040
rect -1162 944 -1128 968
rect -1162 861 -1128 896
rect -704 1434 -670 1469
rect -704 1362 -670 1386
rect -704 1290 -670 1318
rect -704 1218 -670 1250
rect -704 1148 -670 1182
rect -704 1080 -670 1112
rect -704 1012 -670 1040
rect -704 944 -670 968
rect -704 861 -670 896
rect -246 1434 -212 1469
rect -246 1362 -212 1386
rect -246 1290 -212 1318
rect -246 1218 -212 1250
rect -246 1148 -212 1182
rect -246 1080 -212 1112
rect -246 1012 -212 1040
rect -246 944 -212 968
rect -246 861 -212 896
rect 212 1434 246 1469
rect 212 1362 246 1386
rect 212 1290 246 1318
rect 212 1218 246 1250
rect 212 1148 246 1182
rect 212 1080 246 1112
rect 212 1012 246 1040
rect 212 944 246 968
rect 212 861 246 896
rect 670 1434 704 1469
rect 670 1362 704 1386
rect 670 1290 704 1318
rect 670 1218 704 1250
rect 670 1148 704 1182
rect 670 1080 704 1112
rect 670 1012 704 1040
rect 670 944 704 968
rect 670 861 704 896
rect 1128 1434 1162 1469
rect 1128 1362 1162 1386
rect 1128 1290 1162 1318
rect 1128 1218 1162 1250
rect 1128 1148 1162 1182
rect 1128 1080 1162 1112
rect 1128 1012 1162 1040
rect 1128 944 1162 968
rect 1128 861 1162 896
rect -1116 793 -1077 827
rect -1035 793 -1005 827
rect -967 793 -933 827
rect -899 793 -865 827
rect -827 793 -797 827
rect -755 793 -716 827
rect -658 793 -619 827
rect -577 793 -547 827
rect -509 793 -475 827
rect -441 793 -407 827
rect -369 793 -339 827
rect -297 793 -258 827
rect -200 793 -161 827
rect -119 793 -89 827
rect -51 793 -17 827
rect 17 793 51 827
rect 89 793 119 827
rect 161 793 200 827
rect 258 793 297 827
rect 339 793 369 827
rect 407 793 441 827
rect 475 793 509 827
rect 547 793 577 827
rect 619 793 658 827
rect 716 793 755 827
rect 797 793 827 827
rect 865 793 899 827
rect 933 793 967 827
rect 1005 793 1035 827
rect 1077 793 1116 827
rect -1162 678 -1128 713
rect -1162 606 -1128 630
rect -1162 534 -1128 562
rect -1162 462 -1128 494
rect -1162 392 -1128 426
rect -1162 324 -1128 356
rect -1162 256 -1128 284
rect -1162 188 -1128 212
rect -1162 105 -1128 140
rect -704 678 -670 713
rect -704 606 -670 630
rect -704 534 -670 562
rect -704 462 -670 494
rect -704 392 -670 426
rect -704 324 -670 356
rect -704 256 -670 284
rect -704 188 -670 212
rect -704 105 -670 140
rect -246 678 -212 713
rect -246 606 -212 630
rect -246 534 -212 562
rect -246 462 -212 494
rect -246 392 -212 426
rect -246 324 -212 356
rect -246 256 -212 284
rect -246 188 -212 212
rect -246 105 -212 140
rect 212 678 246 713
rect 212 606 246 630
rect 212 534 246 562
rect 212 462 246 494
rect 212 392 246 426
rect 212 324 246 356
rect 212 256 246 284
rect 212 188 246 212
rect 212 105 246 140
rect 670 678 704 713
rect 670 606 704 630
rect 670 534 704 562
rect 670 462 704 494
rect 670 392 704 426
rect 670 324 704 356
rect 670 256 704 284
rect 670 188 704 212
rect 670 105 704 140
rect 1128 678 1162 713
rect 1128 606 1162 630
rect 1128 534 1162 562
rect 1128 462 1162 494
rect 1128 392 1162 426
rect 1128 324 1162 356
rect 1128 256 1162 284
rect 1128 188 1162 212
rect 1128 105 1162 140
rect -1116 37 -1077 71
rect -1035 37 -1005 71
rect -967 37 -933 71
rect -899 37 -865 71
rect -827 37 -797 71
rect -755 37 -716 71
rect -658 37 -619 71
rect -577 37 -547 71
rect -509 37 -475 71
rect -441 37 -407 71
rect -369 37 -339 71
rect -297 37 -258 71
rect -200 37 -161 71
rect -119 37 -89 71
rect -51 37 -17 71
rect 17 37 51 71
rect 89 37 119 71
rect 161 37 200 71
rect 258 37 297 71
rect 339 37 369 71
rect 407 37 441 71
rect 475 37 509 71
rect 547 37 577 71
rect 619 37 658 71
rect 716 37 755 71
rect 797 37 827 71
rect 865 37 899 71
rect 933 37 967 71
rect 1005 37 1035 71
rect 1077 37 1116 71
rect -1162 -78 -1128 -43
rect -1162 -150 -1128 -126
rect -1162 -222 -1128 -194
rect -1162 -294 -1128 -262
rect -1162 -364 -1128 -330
rect -1162 -432 -1128 -400
rect -1162 -500 -1128 -472
rect -1162 -568 -1128 -544
rect -1162 -651 -1128 -616
rect -704 -78 -670 -43
rect -704 -150 -670 -126
rect -704 -222 -670 -194
rect -704 -294 -670 -262
rect -704 -364 -670 -330
rect -704 -432 -670 -400
rect -704 -500 -670 -472
rect -704 -568 -670 -544
rect -704 -651 -670 -616
rect -246 -78 -212 -43
rect -246 -150 -212 -126
rect -246 -222 -212 -194
rect -246 -294 -212 -262
rect -246 -364 -212 -330
rect -246 -432 -212 -400
rect -246 -500 -212 -472
rect -246 -568 -212 -544
rect -246 -651 -212 -616
rect 212 -78 246 -43
rect 212 -150 246 -126
rect 212 -222 246 -194
rect 212 -294 246 -262
rect 212 -364 246 -330
rect 212 -432 246 -400
rect 212 -500 246 -472
rect 212 -568 246 -544
rect 212 -651 246 -616
rect 670 -78 704 -43
rect 670 -150 704 -126
rect 670 -222 704 -194
rect 670 -294 704 -262
rect 670 -364 704 -330
rect 670 -432 704 -400
rect 670 -500 704 -472
rect 670 -568 704 -544
rect 670 -651 704 -616
rect 1128 -78 1162 -43
rect 1128 -150 1162 -126
rect 1128 -222 1162 -194
rect 1128 -294 1162 -262
rect 1128 -364 1162 -330
rect 1128 -432 1162 -400
rect 1128 -500 1162 -472
rect 1128 -568 1162 -544
rect 1128 -651 1162 -616
rect -1116 -719 -1077 -685
rect -1035 -719 -1005 -685
rect -967 -719 -933 -685
rect -899 -719 -865 -685
rect -827 -719 -797 -685
rect -755 -719 -716 -685
rect -658 -719 -619 -685
rect -577 -719 -547 -685
rect -509 -719 -475 -685
rect -441 -719 -407 -685
rect -369 -719 -339 -685
rect -297 -719 -258 -685
rect -200 -719 -161 -685
rect -119 -719 -89 -685
rect -51 -719 -17 -685
rect 17 -719 51 -685
rect 89 -719 119 -685
rect 161 -719 200 -685
rect 258 -719 297 -685
rect 339 -719 369 -685
rect 407 -719 441 -685
rect 475 -719 509 -685
rect 547 -719 577 -685
rect 619 -719 658 -685
rect 716 -719 755 -685
rect 797 -719 827 -685
rect 865 -719 899 -685
rect 933 -719 967 -685
rect 1005 -719 1035 -685
rect 1077 -719 1116 -685
rect -1162 -834 -1128 -799
rect -1162 -906 -1128 -882
rect -1162 -978 -1128 -950
rect -1162 -1050 -1128 -1018
rect -1162 -1120 -1128 -1086
rect -1162 -1188 -1128 -1156
rect -1162 -1256 -1128 -1228
rect -1162 -1324 -1128 -1300
rect -1162 -1407 -1128 -1372
rect -704 -834 -670 -799
rect -704 -906 -670 -882
rect -704 -978 -670 -950
rect -704 -1050 -670 -1018
rect -704 -1120 -670 -1086
rect -704 -1188 -670 -1156
rect -704 -1256 -670 -1228
rect -704 -1324 -670 -1300
rect -704 -1407 -670 -1372
rect -246 -834 -212 -799
rect -246 -906 -212 -882
rect -246 -978 -212 -950
rect -246 -1050 -212 -1018
rect -246 -1120 -212 -1086
rect -246 -1188 -212 -1156
rect -246 -1256 -212 -1228
rect -246 -1324 -212 -1300
rect -246 -1407 -212 -1372
rect 212 -834 246 -799
rect 212 -906 246 -882
rect 212 -978 246 -950
rect 212 -1050 246 -1018
rect 212 -1120 246 -1086
rect 212 -1188 246 -1156
rect 212 -1256 246 -1228
rect 212 -1324 246 -1300
rect 212 -1407 246 -1372
rect 670 -834 704 -799
rect 670 -906 704 -882
rect 670 -978 704 -950
rect 670 -1050 704 -1018
rect 670 -1120 704 -1086
rect 670 -1188 704 -1156
rect 670 -1256 704 -1228
rect 670 -1324 704 -1300
rect 670 -1407 704 -1372
rect 1128 -834 1162 -799
rect 1128 -906 1162 -882
rect 1128 -978 1162 -950
rect 1128 -1050 1162 -1018
rect 1128 -1120 1162 -1086
rect 1128 -1188 1162 -1156
rect 1128 -1256 1162 -1228
rect 1128 -1324 1162 -1300
rect 1128 -1407 1162 -1372
rect -1116 -1475 -1077 -1441
rect -1035 -1475 -1005 -1441
rect -967 -1475 -933 -1441
rect -899 -1475 -865 -1441
rect -827 -1475 -797 -1441
rect -755 -1475 -716 -1441
rect -658 -1475 -619 -1441
rect -577 -1475 -547 -1441
rect -509 -1475 -475 -1441
rect -441 -1475 -407 -1441
rect -369 -1475 -339 -1441
rect -297 -1475 -258 -1441
rect -200 -1475 -161 -1441
rect -119 -1475 -89 -1441
rect -51 -1475 -17 -1441
rect 17 -1475 51 -1441
rect 89 -1475 119 -1441
rect 161 -1475 200 -1441
rect 258 -1475 297 -1441
rect 339 -1475 369 -1441
rect 407 -1475 441 -1441
rect 475 -1475 509 -1441
rect 547 -1475 577 -1441
rect 619 -1475 658 -1441
rect 716 -1475 755 -1441
rect 797 -1475 827 -1441
rect 865 -1475 899 -1441
rect 933 -1475 967 -1441
rect 1005 -1475 1035 -1441
rect 1077 -1475 1116 -1441
rect 1242 -1543 1276 1543
rect -1276 -1577 -1173 -1543
rect -1139 -1577 -1105 -1543
rect -1071 -1577 -1037 -1543
rect -1003 -1577 -969 -1543
rect -935 -1577 -901 -1543
rect -867 -1577 -833 -1543
rect -799 -1577 -765 -1543
rect -731 -1577 -697 -1543
rect -663 -1577 -629 -1543
rect -595 -1577 -561 -1543
rect -527 -1577 -493 -1543
rect -459 -1577 -425 -1543
rect -391 -1577 -357 -1543
rect -323 -1577 -289 -1543
rect -255 -1577 -221 -1543
rect -187 -1577 -153 -1543
rect -119 -1577 -85 -1543
rect -51 -1577 -17 -1543
rect 17 -1577 51 -1543
rect 85 -1577 119 -1543
rect 153 -1577 187 -1543
rect 221 -1577 255 -1543
rect 289 -1577 323 -1543
rect 357 -1577 391 -1543
rect 425 -1577 459 -1543
rect 493 -1577 527 -1543
rect 561 -1577 595 -1543
rect 629 -1577 663 -1543
rect 697 -1577 731 -1543
rect 765 -1577 799 -1543
rect 833 -1577 867 -1543
rect 901 -1577 935 -1543
rect 969 -1577 1003 -1543
rect 1037 -1577 1071 -1543
rect 1105 -1577 1139 -1543
rect 1173 -1577 1276 -1543
<< viali >>
rect -1162 1420 -1128 1434
rect -1162 1400 -1128 1420
rect -1162 1352 -1128 1362
rect -1162 1328 -1128 1352
rect -1162 1284 -1128 1290
rect -1162 1256 -1128 1284
rect -1162 1216 -1128 1218
rect -1162 1184 -1128 1216
rect -1162 1114 -1128 1146
rect -1162 1112 -1128 1114
rect -1162 1046 -1128 1074
rect -1162 1040 -1128 1046
rect -1162 978 -1128 1002
rect -1162 968 -1128 978
rect -1162 910 -1128 930
rect -1162 896 -1128 910
rect -704 1420 -670 1434
rect -704 1400 -670 1420
rect -704 1352 -670 1362
rect -704 1328 -670 1352
rect -704 1284 -670 1290
rect -704 1256 -670 1284
rect -704 1216 -670 1218
rect -704 1184 -670 1216
rect -704 1114 -670 1146
rect -704 1112 -670 1114
rect -704 1046 -670 1074
rect -704 1040 -670 1046
rect -704 978 -670 1002
rect -704 968 -670 978
rect -704 910 -670 930
rect -704 896 -670 910
rect -246 1420 -212 1434
rect -246 1400 -212 1420
rect -246 1352 -212 1362
rect -246 1328 -212 1352
rect -246 1284 -212 1290
rect -246 1256 -212 1284
rect -246 1216 -212 1218
rect -246 1184 -212 1216
rect -246 1114 -212 1146
rect -246 1112 -212 1114
rect -246 1046 -212 1074
rect -246 1040 -212 1046
rect -246 978 -212 1002
rect -246 968 -212 978
rect -246 910 -212 930
rect -246 896 -212 910
rect 212 1420 246 1434
rect 212 1400 246 1420
rect 212 1352 246 1362
rect 212 1328 246 1352
rect 212 1284 246 1290
rect 212 1256 246 1284
rect 212 1216 246 1218
rect 212 1184 246 1216
rect 212 1114 246 1146
rect 212 1112 246 1114
rect 212 1046 246 1074
rect 212 1040 246 1046
rect 212 978 246 1002
rect 212 968 246 978
rect 212 910 246 930
rect 212 896 246 910
rect 670 1420 704 1434
rect 670 1400 704 1420
rect 670 1352 704 1362
rect 670 1328 704 1352
rect 670 1284 704 1290
rect 670 1256 704 1284
rect 670 1216 704 1218
rect 670 1184 704 1216
rect 670 1114 704 1146
rect 670 1112 704 1114
rect 670 1046 704 1074
rect 670 1040 704 1046
rect 670 978 704 1002
rect 670 968 704 978
rect 670 910 704 930
rect 670 896 704 910
rect 1128 1420 1162 1434
rect 1128 1400 1162 1420
rect 1128 1352 1162 1362
rect 1128 1328 1162 1352
rect 1128 1284 1162 1290
rect 1128 1256 1162 1284
rect 1128 1216 1162 1218
rect 1128 1184 1162 1216
rect 1128 1114 1162 1146
rect 1128 1112 1162 1114
rect 1128 1046 1162 1074
rect 1128 1040 1162 1046
rect 1128 978 1162 1002
rect 1128 968 1162 978
rect 1128 910 1162 930
rect 1128 896 1162 910
rect -1077 793 -1069 827
rect -1069 793 -1043 827
rect -1005 793 -1001 827
rect -1001 793 -971 827
rect -933 793 -899 827
rect -861 793 -831 827
rect -831 793 -827 827
rect -789 793 -763 827
rect -763 793 -755 827
rect -619 793 -611 827
rect -611 793 -585 827
rect -547 793 -543 827
rect -543 793 -513 827
rect -475 793 -441 827
rect -403 793 -373 827
rect -373 793 -369 827
rect -331 793 -305 827
rect -305 793 -297 827
rect -161 793 -153 827
rect -153 793 -127 827
rect -89 793 -85 827
rect -85 793 -55 827
rect -17 793 17 827
rect 55 793 85 827
rect 85 793 89 827
rect 127 793 153 827
rect 153 793 161 827
rect 297 793 305 827
rect 305 793 331 827
rect 369 793 373 827
rect 373 793 403 827
rect 441 793 475 827
rect 513 793 543 827
rect 543 793 547 827
rect 585 793 611 827
rect 611 793 619 827
rect 755 793 763 827
rect 763 793 789 827
rect 827 793 831 827
rect 831 793 861 827
rect 899 793 933 827
rect 971 793 1001 827
rect 1001 793 1005 827
rect 1043 793 1069 827
rect 1069 793 1077 827
rect -1162 664 -1128 678
rect -1162 644 -1128 664
rect -1162 596 -1128 606
rect -1162 572 -1128 596
rect -1162 528 -1128 534
rect -1162 500 -1128 528
rect -1162 460 -1128 462
rect -1162 428 -1128 460
rect -1162 358 -1128 390
rect -1162 356 -1128 358
rect -1162 290 -1128 318
rect -1162 284 -1128 290
rect -1162 222 -1128 246
rect -1162 212 -1128 222
rect -1162 154 -1128 174
rect -1162 140 -1128 154
rect -704 664 -670 678
rect -704 644 -670 664
rect -704 596 -670 606
rect -704 572 -670 596
rect -704 528 -670 534
rect -704 500 -670 528
rect -704 460 -670 462
rect -704 428 -670 460
rect -704 358 -670 390
rect -704 356 -670 358
rect -704 290 -670 318
rect -704 284 -670 290
rect -704 222 -670 246
rect -704 212 -670 222
rect -704 154 -670 174
rect -704 140 -670 154
rect -246 664 -212 678
rect -246 644 -212 664
rect -246 596 -212 606
rect -246 572 -212 596
rect -246 528 -212 534
rect -246 500 -212 528
rect -246 460 -212 462
rect -246 428 -212 460
rect -246 358 -212 390
rect -246 356 -212 358
rect -246 290 -212 318
rect -246 284 -212 290
rect -246 222 -212 246
rect -246 212 -212 222
rect -246 154 -212 174
rect -246 140 -212 154
rect 212 664 246 678
rect 212 644 246 664
rect 212 596 246 606
rect 212 572 246 596
rect 212 528 246 534
rect 212 500 246 528
rect 212 460 246 462
rect 212 428 246 460
rect 212 358 246 390
rect 212 356 246 358
rect 212 290 246 318
rect 212 284 246 290
rect 212 222 246 246
rect 212 212 246 222
rect 212 154 246 174
rect 212 140 246 154
rect 670 664 704 678
rect 670 644 704 664
rect 670 596 704 606
rect 670 572 704 596
rect 670 528 704 534
rect 670 500 704 528
rect 670 460 704 462
rect 670 428 704 460
rect 670 358 704 390
rect 670 356 704 358
rect 670 290 704 318
rect 670 284 704 290
rect 670 222 704 246
rect 670 212 704 222
rect 670 154 704 174
rect 670 140 704 154
rect 1128 664 1162 678
rect 1128 644 1162 664
rect 1128 596 1162 606
rect 1128 572 1162 596
rect 1128 528 1162 534
rect 1128 500 1162 528
rect 1128 460 1162 462
rect 1128 428 1162 460
rect 1128 358 1162 390
rect 1128 356 1162 358
rect 1128 290 1162 318
rect 1128 284 1162 290
rect 1128 222 1162 246
rect 1128 212 1162 222
rect 1128 154 1162 174
rect 1128 140 1162 154
rect -1077 37 -1069 71
rect -1069 37 -1043 71
rect -1005 37 -1001 71
rect -1001 37 -971 71
rect -933 37 -899 71
rect -861 37 -831 71
rect -831 37 -827 71
rect -789 37 -763 71
rect -763 37 -755 71
rect -619 37 -611 71
rect -611 37 -585 71
rect -547 37 -543 71
rect -543 37 -513 71
rect -475 37 -441 71
rect -403 37 -373 71
rect -373 37 -369 71
rect -331 37 -305 71
rect -305 37 -297 71
rect -161 37 -153 71
rect -153 37 -127 71
rect -89 37 -85 71
rect -85 37 -55 71
rect -17 37 17 71
rect 55 37 85 71
rect 85 37 89 71
rect 127 37 153 71
rect 153 37 161 71
rect 297 37 305 71
rect 305 37 331 71
rect 369 37 373 71
rect 373 37 403 71
rect 441 37 475 71
rect 513 37 543 71
rect 543 37 547 71
rect 585 37 611 71
rect 611 37 619 71
rect 755 37 763 71
rect 763 37 789 71
rect 827 37 831 71
rect 831 37 861 71
rect 899 37 933 71
rect 971 37 1001 71
rect 1001 37 1005 71
rect 1043 37 1069 71
rect 1069 37 1077 71
rect -1162 -92 -1128 -78
rect -1162 -112 -1128 -92
rect -1162 -160 -1128 -150
rect -1162 -184 -1128 -160
rect -1162 -228 -1128 -222
rect -1162 -256 -1128 -228
rect -1162 -296 -1128 -294
rect -1162 -328 -1128 -296
rect -1162 -398 -1128 -366
rect -1162 -400 -1128 -398
rect -1162 -466 -1128 -438
rect -1162 -472 -1128 -466
rect -1162 -534 -1128 -510
rect -1162 -544 -1128 -534
rect -1162 -602 -1128 -582
rect -1162 -616 -1128 -602
rect -704 -92 -670 -78
rect -704 -112 -670 -92
rect -704 -160 -670 -150
rect -704 -184 -670 -160
rect -704 -228 -670 -222
rect -704 -256 -670 -228
rect -704 -296 -670 -294
rect -704 -328 -670 -296
rect -704 -398 -670 -366
rect -704 -400 -670 -398
rect -704 -466 -670 -438
rect -704 -472 -670 -466
rect -704 -534 -670 -510
rect -704 -544 -670 -534
rect -704 -602 -670 -582
rect -704 -616 -670 -602
rect -246 -92 -212 -78
rect -246 -112 -212 -92
rect -246 -160 -212 -150
rect -246 -184 -212 -160
rect -246 -228 -212 -222
rect -246 -256 -212 -228
rect -246 -296 -212 -294
rect -246 -328 -212 -296
rect -246 -398 -212 -366
rect -246 -400 -212 -398
rect -246 -466 -212 -438
rect -246 -472 -212 -466
rect -246 -534 -212 -510
rect -246 -544 -212 -534
rect -246 -602 -212 -582
rect -246 -616 -212 -602
rect 212 -92 246 -78
rect 212 -112 246 -92
rect 212 -160 246 -150
rect 212 -184 246 -160
rect 212 -228 246 -222
rect 212 -256 246 -228
rect 212 -296 246 -294
rect 212 -328 246 -296
rect 212 -398 246 -366
rect 212 -400 246 -398
rect 212 -466 246 -438
rect 212 -472 246 -466
rect 212 -534 246 -510
rect 212 -544 246 -534
rect 212 -602 246 -582
rect 212 -616 246 -602
rect 670 -92 704 -78
rect 670 -112 704 -92
rect 670 -160 704 -150
rect 670 -184 704 -160
rect 670 -228 704 -222
rect 670 -256 704 -228
rect 670 -296 704 -294
rect 670 -328 704 -296
rect 670 -398 704 -366
rect 670 -400 704 -398
rect 670 -466 704 -438
rect 670 -472 704 -466
rect 670 -534 704 -510
rect 670 -544 704 -534
rect 670 -602 704 -582
rect 670 -616 704 -602
rect 1128 -92 1162 -78
rect 1128 -112 1162 -92
rect 1128 -160 1162 -150
rect 1128 -184 1162 -160
rect 1128 -228 1162 -222
rect 1128 -256 1162 -228
rect 1128 -296 1162 -294
rect 1128 -328 1162 -296
rect 1128 -398 1162 -366
rect 1128 -400 1162 -398
rect 1128 -466 1162 -438
rect 1128 -472 1162 -466
rect 1128 -534 1162 -510
rect 1128 -544 1162 -534
rect 1128 -602 1162 -582
rect 1128 -616 1162 -602
rect -1077 -719 -1069 -685
rect -1069 -719 -1043 -685
rect -1005 -719 -1001 -685
rect -1001 -719 -971 -685
rect -933 -719 -899 -685
rect -861 -719 -831 -685
rect -831 -719 -827 -685
rect -789 -719 -763 -685
rect -763 -719 -755 -685
rect -619 -719 -611 -685
rect -611 -719 -585 -685
rect -547 -719 -543 -685
rect -543 -719 -513 -685
rect -475 -719 -441 -685
rect -403 -719 -373 -685
rect -373 -719 -369 -685
rect -331 -719 -305 -685
rect -305 -719 -297 -685
rect -161 -719 -153 -685
rect -153 -719 -127 -685
rect -89 -719 -85 -685
rect -85 -719 -55 -685
rect -17 -719 17 -685
rect 55 -719 85 -685
rect 85 -719 89 -685
rect 127 -719 153 -685
rect 153 -719 161 -685
rect 297 -719 305 -685
rect 305 -719 331 -685
rect 369 -719 373 -685
rect 373 -719 403 -685
rect 441 -719 475 -685
rect 513 -719 543 -685
rect 543 -719 547 -685
rect 585 -719 611 -685
rect 611 -719 619 -685
rect 755 -719 763 -685
rect 763 -719 789 -685
rect 827 -719 831 -685
rect 831 -719 861 -685
rect 899 -719 933 -685
rect 971 -719 1001 -685
rect 1001 -719 1005 -685
rect 1043 -719 1069 -685
rect 1069 -719 1077 -685
rect -1162 -848 -1128 -834
rect -1162 -868 -1128 -848
rect -1162 -916 -1128 -906
rect -1162 -940 -1128 -916
rect -1162 -984 -1128 -978
rect -1162 -1012 -1128 -984
rect -1162 -1052 -1128 -1050
rect -1162 -1084 -1128 -1052
rect -1162 -1154 -1128 -1122
rect -1162 -1156 -1128 -1154
rect -1162 -1222 -1128 -1194
rect -1162 -1228 -1128 -1222
rect -1162 -1290 -1128 -1266
rect -1162 -1300 -1128 -1290
rect -1162 -1358 -1128 -1338
rect -1162 -1372 -1128 -1358
rect -704 -848 -670 -834
rect -704 -868 -670 -848
rect -704 -916 -670 -906
rect -704 -940 -670 -916
rect -704 -984 -670 -978
rect -704 -1012 -670 -984
rect -704 -1052 -670 -1050
rect -704 -1084 -670 -1052
rect -704 -1154 -670 -1122
rect -704 -1156 -670 -1154
rect -704 -1222 -670 -1194
rect -704 -1228 -670 -1222
rect -704 -1290 -670 -1266
rect -704 -1300 -670 -1290
rect -704 -1358 -670 -1338
rect -704 -1372 -670 -1358
rect -246 -848 -212 -834
rect -246 -868 -212 -848
rect -246 -916 -212 -906
rect -246 -940 -212 -916
rect -246 -984 -212 -978
rect -246 -1012 -212 -984
rect -246 -1052 -212 -1050
rect -246 -1084 -212 -1052
rect -246 -1154 -212 -1122
rect -246 -1156 -212 -1154
rect -246 -1222 -212 -1194
rect -246 -1228 -212 -1222
rect -246 -1290 -212 -1266
rect -246 -1300 -212 -1290
rect -246 -1358 -212 -1338
rect -246 -1372 -212 -1358
rect 212 -848 246 -834
rect 212 -868 246 -848
rect 212 -916 246 -906
rect 212 -940 246 -916
rect 212 -984 246 -978
rect 212 -1012 246 -984
rect 212 -1052 246 -1050
rect 212 -1084 246 -1052
rect 212 -1154 246 -1122
rect 212 -1156 246 -1154
rect 212 -1222 246 -1194
rect 212 -1228 246 -1222
rect 212 -1290 246 -1266
rect 212 -1300 246 -1290
rect 212 -1358 246 -1338
rect 212 -1372 246 -1358
rect 670 -848 704 -834
rect 670 -868 704 -848
rect 670 -916 704 -906
rect 670 -940 704 -916
rect 670 -984 704 -978
rect 670 -1012 704 -984
rect 670 -1052 704 -1050
rect 670 -1084 704 -1052
rect 670 -1154 704 -1122
rect 670 -1156 704 -1154
rect 670 -1222 704 -1194
rect 670 -1228 704 -1222
rect 670 -1290 704 -1266
rect 670 -1300 704 -1290
rect 670 -1358 704 -1338
rect 670 -1372 704 -1358
rect 1128 -848 1162 -834
rect 1128 -868 1162 -848
rect 1128 -916 1162 -906
rect 1128 -940 1162 -916
rect 1128 -984 1162 -978
rect 1128 -1012 1162 -984
rect 1128 -1052 1162 -1050
rect 1128 -1084 1162 -1052
rect 1128 -1154 1162 -1122
rect 1128 -1156 1162 -1154
rect 1128 -1222 1162 -1194
rect 1128 -1228 1162 -1222
rect 1128 -1290 1162 -1266
rect 1128 -1300 1162 -1290
rect 1128 -1358 1162 -1338
rect 1128 -1372 1162 -1358
rect -1077 -1475 -1069 -1441
rect -1069 -1475 -1043 -1441
rect -1005 -1475 -1001 -1441
rect -1001 -1475 -971 -1441
rect -933 -1475 -899 -1441
rect -861 -1475 -831 -1441
rect -831 -1475 -827 -1441
rect -789 -1475 -763 -1441
rect -763 -1475 -755 -1441
rect -619 -1475 -611 -1441
rect -611 -1475 -585 -1441
rect -547 -1475 -543 -1441
rect -543 -1475 -513 -1441
rect -475 -1475 -441 -1441
rect -403 -1475 -373 -1441
rect -373 -1475 -369 -1441
rect -331 -1475 -305 -1441
rect -305 -1475 -297 -1441
rect -161 -1475 -153 -1441
rect -153 -1475 -127 -1441
rect -89 -1475 -85 -1441
rect -85 -1475 -55 -1441
rect -17 -1475 17 -1441
rect 55 -1475 85 -1441
rect 85 -1475 89 -1441
rect 127 -1475 153 -1441
rect 153 -1475 161 -1441
rect 297 -1475 305 -1441
rect 305 -1475 331 -1441
rect 369 -1475 373 -1441
rect 373 -1475 403 -1441
rect 441 -1475 475 -1441
rect 513 -1475 543 -1441
rect 543 -1475 547 -1441
rect 585 -1475 611 -1441
rect 611 -1475 619 -1441
rect 755 -1475 763 -1441
rect 763 -1475 789 -1441
rect 827 -1475 831 -1441
rect 831 -1475 861 -1441
rect 899 -1475 933 -1441
rect 971 -1475 1001 -1441
rect 1001 -1475 1005 -1441
rect 1043 -1475 1069 -1441
rect 1069 -1475 1077 -1441
<< metal1 >>
rect -1168 1434 -1122 1465
rect -1168 1400 -1162 1434
rect -1128 1400 -1122 1434
rect -1168 1362 -1122 1400
rect -1168 1328 -1162 1362
rect -1128 1328 -1122 1362
rect -1168 1290 -1122 1328
rect -1168 1256 -1162 1290
rect -1128 1256 -1122 1290
rect -1168 1218 -1122 1256
rect -1168 1184 -1162 1218
rect -1128 1184 -1122 1218
rect -1168 1146 -1122 1184
rect -1168 1112 -1162 1146
rect -1128 1112 -1122 1146
rect -1168 1074 -1122 1112
rect -1168 1040 -1162 1074
rect -1128 1040 -1122 1074
rect -1168 1002 -1122 1040
rect -1168 968 -1162 1002
rect -1128 968 -1122 1002
rect -1168 930 -1122 968
rect -1168 896 -1162 930
rect -1128 896 -1122 930
rect -1168 865 -1122 896
rect -710 1434 -664 1465
rect -710 1400 -704 1434
rect -670 1400 -664 1434
rect -710 1362 -664 1400
rect -710 1328 -704 1362
rect -670 1328 -664 1362
rect -710 1290 -664 1328
rect -710 1256 -704 1290
rect -670 1256 -664 1290
rect -710 1218 -664 1256
rect -710 1184 -704 1218
rect -670 1184 -664 1218
rect -710 1146 -664 1184
rect -710 1112 -704 1146
rect -670 1112 -664 1146
rect -710 1074 -664 1112
rect -710 1040 -704 1074
rect -670 1040 -664 1074
rect -710 1002 -664 1040
rect -710 968 -704 1002
rect -670 968 -664 1002
rect -710 930 -664 968
rect -710 896 -704 930
rect -670 896 -664 930
rect -710 865 -664 896
rect -252 1434 -206 1465
rect -252 1400 -246 1434
rect -212 1400 -206 1434
rect -252 1362 -206 1400
rect -252 1328 -246 1362
rect -212 1328 -206 1362
rect -252 1290 -206 1328
rect -252 1256 -246 1290
rect -212 1256 -206 1290
rect -252 1218 -206 1256
rect -252 1184 -246 1218
rect -212 1184 -206 1218
rect -252 1146 -206 1184
rect -252 1112 -246 1146
rect -212 1112 -206 1146
rect -252 1074 -206 1112
rect -252 1040 -246 1074
rect -212 1040 -206 1074
rect -252 1002 -206 1040
rect -252 968 -246 1002
rect -212 968 -206 1002
rect -252 930 -206 968
rect -252 896 -246 930
rect -212 896 -206 930
rect -252 865 -206 896
rect 206 1434 252 1465
rect 206 1400 212 1434
rect 246 1400 252 1434
rect 206 1362 252 1400
rect 206 1328 212 1362
rect 246 1328 252 1362
rect 206 1290 252 1328
rect 206 1256 212 1290
rect 246 1256 252 1290
rect 206 1218 252 1256
rect 206 1184 212 1218
rect 246 1184 252 1218
rect 206 1146 252 1184
rect 206 1112 212 1146
rect 246 1112 252 1146
rect 206 1074 252 1112
rect 206 1040 212 1074
rect 246 1040 252 1074
rect 206 1002 252 1040
rect 206 968 212 1002
rect 246 968 252 1002
rect 206 930 252 968
rect 206 896 212 930
rect 246 896 252 930
rect 206 865 252 896
rect 664 1434 710 1465
rect 664 1400 670 1434
rect 704 1400 710 1434
rect 664 1362 710 1400
rect 664 1328 670 1362
rect 704 1328 710 1362
rect 664 1290 710 1328
rect 664 1256 670 1290
rect 704 1256 710 1290
rect 664 1218 710 1256
rect 664 1184 670 1218
rect 704 1184 710 1218
rect 664 1146 710 1184
rect 664 1112 670 1146
rect 704 1112 710 1146
rect 664 1074 710 1112
rect 664 1040 670 1074
rect 704 1040 710 1074
rect 664 1002 710 1040
rect 664 968 670 1002
rect 704 968 710 1002
rect 664 930 710 968
rect 664 896 670 930
rect 704 896 710 930
rect 664 865 710 896
rect 1122 1434 1168 1465
rect 1122 1400 1128 1434
rect 1162 1400 1168 1434
rect 1122 1362 1168 1400
rect 1122 1328 1128 1362
rect 1162 1328 1168 1362
rect 1122 1290 1168 1328
rect 1122 1256 1128 1290
rect 1162 1256 1168 1290
rect 1122 1218 1168 1256
rect 1122 1184 1128 1218
rect 1162 1184 1168 1218
rect 1122 1146 1168 1184
rect 1122 1112 1128 1146
rect 1162 1112 1168 1146
rect 1122 1074 1168 1112
rect 1122 1040 1128 1074
rect 1162 1040 1168 1074
rect 1122 1002 1168 1040
rect 1122 968 1128 1002
rect 1162 968 1168 1002
rect 1122 930 1168 968
rect 1122 896 1128 930
rect 1162 896 1168 930
rect 1122 865 1168 896
rect -1112 827 -720 833
rect -1112 793 -1077 827
rect -1043 793 -1005 827
rect -971 793 -933 827
rect -899 793 -861 827
rect -827 793 -789 827
rect -755 793 -720 827
rect -1112 787 -720 793
rect -654 827 -262 833
rect -654 793 -619 827
rect -585 793 -547 827
rect -513 793 -475 827
rect -441 793 -403 827
rect -369 793 -331 827
rect -297 793 -262 827
rect -654 787 -262 793
rect -196 827 196 833
rect -196 793 -161 827
rect -127 793 -89 827
rect -55 793 -17 827
rect 17 793 55 827
rect 89 793 127 827
rect 161 793 196 827
rect -196 787 196 793
rect 262 827 654 833
rect 262 793 297 827
rect 331 793 369 827
rect 403 793 441 827
rect 475 793 513 827
rect 547 793 585 827
rect 619 793 654 827
rect 262 787 654 793
rect 720 827 1112 833
rect 720 793 755 827
rect 789 793 827 827
rect 861 793 899 827
rect 933 793 971 827
rect 1005 793 1043 827
rect 1077 793 1112 827
rect 720 787 1112 793
rect -1168 678 -1122 709
rect -1168 644 -1162 678
rect -1128 644 -1122 678
rect -1168 606 -1122 644
rect -1168 572 -1162 606
rect -1128 572 -1122 606
rect -1168 534 -1122 572
rect -1168 500 -1162 534
rect -1128 500 -1122 534
rect -1168 462 -1122 500
rect -1168 428 -1162 462
rect -1128 428 -1122 462
rect -1168 390 -1122 428
rect -1168 356 -1162 390
rect -1128 356 -1122 390
rect -1168 318 -1122 356
rect -1168 284 -1162 318
rect -1128 284 -1122 318
rect -1168 246 -1122 284
rect -1168 212 -1162 246
rect -1128 212 -1122 246
rect -1168 174 -1122 212
rect -1168 140 -1162 174
rect -1128 140 -1122 174
rect -1168 109 -1122 140
rect -710 678 -664 709
rect -710 644 -704 678
rect -670 644 -664 678
rect -710 606 -664 644
rect -710 572 -704 606
rect -670 572 -664 606
rect -710 534 -664 572
rect -710 500 -704 534
rect -670 500 -664 534
rect -710 462 -664 500
rect -710 428 -704 462
rect -670 428 -664 462
rect -710 390 -664 428
rect -710 356 -704 390
rect -670 356 -664 390
rect -710 318 -664 356
rect -710 284 -704 318
rect -670 284 -664 318
rect -710 246 -664 284
rect -710 212 -704 246
rect -670 212 -664 246
rect -710 174 -664 212
rect -710 140 -704 174
rect -670 140 -664 174
rect -710 109 -664 140
rect -252 678 -206 709
rect -252 644 -246 678
rect -212 644 -206 678
rect -252 606 -206 644
rect -252 572 -246 606
rect -212 572 -206 606
rect -252 534 -206 572
rect -252 500 -246 534
rect -212 500 -206 534
rect -252 462 -206 500
rect -252 428 -246 462
rect -212 428 -206 462
rect -252 390 -206 428
rect -252 356 -246 390
rect -212 356 -206 390
rect -252 318 -206 356
rect -252 284 -246 318
rect -212 284 -206 318
rect -252 246 -206 284
rect -252 212 -246 246
rect -212 212 -206 246
rect -252 174 -206 212
rect -252 140 -246 174
rect -212 140 -206 174
rect -252 109 -206 140
rect 206 678 252 709
rect 206 644 212 678
rect 246 644 252 678
rect 206 606 252 644
rect 206 572 212 606
rect 246 572 252 606
rect 206 534 252 572
rect 206 500 212 534
rect 246 500 252 534
rect 206 462 252 500
rect 206 428 212 462
rect 246 428 252 462
rect 206 390 252 428
rect 206 356 212 390
rect 246 356 252 390
rect 206 318 252 356
rect 206 284 212 318
rect 246 284 252 318
rect 206 246 252 284
rect 206 212 212 246
rect 246 212 252 246
rect 206 174 252 212
rect 206 140 212 174
rect 246 140 252 174
rect 206 109 252 140
rect 664 678 710 709
rect 664 644 670 678
rect 704 644 710 678
rect 664 606 710 644
rect 664 572 670 606
rect 704 572 710 606
rect 664 534 710 572
rect 664 500 670 534
rect 704 500 710 534
rect 664 462 710 500
rect 664 428 670 462
rect 704 428 710 462
rect 664 390 710 428
rect 664 356 670 390
rect 704 356 710 390
rect 664 318 710 356
rect 664 284 670 318
rect 704 284 710 318
rect 664 246 710 284
rect 664 212 670 246
rect 704 212 710 246
rect 664 174 710 212
rect 664 140 670 174
rect 704 140 710 174
rect 664 109 710 140
rect 1122 678 1168 709
rect 1122 644 1128 678
rect 1162 644 1168 678
rect 1122 606 1168 644
rect 1122 572 1128 606
rect 1162 572 1168 606
rect 1122 534 1168 572
rect 1122 500 1128 534
rect 1162 500 1168 534
rect 1122 462 1168 500
rect 1122 428 1128 462
rect 1162 428 1168 462
rect 1122 390 1168 428
rect 1122 356 1128 390
rect 1162 356 1168 390
rect 1122 318 1168 356
rect 1122 284 1128 318
rect 1162 284 1168 318
rect 1122 246 1168 284
rect 1122 212 1128 246
rect 1162 212 1168 246
rect 1122 174 1168 212
rect 1122 140 1128 174
rect 1162 140 1168 174
rect 1122 109 1168 140
rect -1112 71 -720 77
rect -1112 37 -1077 71
rect -1043 37 -1005 71
rect -971 37 -933 71
rect -899 37 -861 71
rect -827 37 -789 71
rect -755 37 -720 71
rect -1112 31 -720 37
rect -654 71 -262 77
rect -654 37 -619 71
rect -585 37 -547 71
rect -513 37 -475 71
rect -441 37 -403 71
rect -369 37 -331 71
rect -297 37 -262 71
rect -654 31 -262 37
rect -196 71 196 77
rect -196 37 -161 71
rect -127 37 -89 71
rect -55 37 -17 71
rect 17 37 55 71
rect 89 37 127 71
rect 161 37 196 71
rect -196 31 196 37
rect 262 71 654 77
rect 262 37 297 71
rect 331 37 369 71
rect 403 37 441 71
rect 475 37 513 71
rect 547 37 585 71
rect 619 37 654 71
rect 262 31 654 37
rect 720 71 1112 77
rect 720 37 755 71
rect 789 37 827 71
rect 861 37 899 71
rect 933 37 971 71
rect 1005 37 1043 71
rect 1077 37 1112 71
rect 720 31 1112 37
rect -1168 -78 -1122 -47
rect -1168 -112 -1162 -78
rect -1128 -112 -1122 -78
rect -1168 -150 -1122 -112
rect -1168 -184 -1162 -150
rect -1128 -184 -1122 -150
rect -1168 -222 -1122 -184
rect -1168 -256 -1162 -222
rect -1128 -256 -1122 -222
rect -1168 -294 -1122 -256
rect -1168 -328 -1162 -294
rect -1128 -328 -1122 -294
rect -1168 -366 -1122 -328
rect -1168 -400 -1162 -366
rect -1128 -400 -1122 -366
rect -1168 -438 -1122 -400
rect -1168 -472 -1162 -438
rect -1128 -472 -1122 -438
rect -1168 -510 -1122 -472
rect -1168 -544 -1162 -510
rect -1128 -544 -1122 -510
rect -1168 -582 -1122 -544
rect -1168 -616 -1162 -582
rect -1128 -616 -1122 -582
rect -1168 -647 -1122 -616
rect -710 -78 -664 -47
rect -710 -112 -704 -78
rect -670 -112 -664 -78
rect -710 -150 -664 -112
rect -710 -184 -704 -150
rect -670 -184 -664 -150
rect -710 -222 -664 -184
rect -710 -256 -704 -222
rect -670 -256 -664 -222
rect -710 -294 -664 -256
rect -710 -328 -704 -294
rect -670 -328 -664 -294
rect -710 -366 -664 -328
rect -710 -400 -704 -366
rect -670 -400 -664 -366
rect -710 -438 -664 -400
rect -710 -472 -704 -438
rect -670 -472 -664 -438
rect -710 -510 -664 -472
rect -710 -544 -704 -510
rect -670 -544 -664 -510
rect -710 -582 -664 -544
rect -710 -616 -704 -582
rect -670 -616 -664 -582
rect -710 -647 -664 -616
rect -252 -78 -206 -47
rect -252 -112 -246 -78
rect -212 -112 -206 -78
rect -252 -150 -206 -112
rect -252 -184 -246 -150
rect -212 -184 -206 -150
rect -252 -222 -206 -184
rect -252 -256 -246 -222
rect -212 -256 -206 -222
rect -252 -294 -206 -256
rect -252 -328 -246 -294
rect -212 -328 -206 -294
rect -252 -366 -206 -328
rect -252 -400 -246 -366
rect -212 -400 -206 -366
rect -252 -438 -206 -400
rect -252 -472 -246 -438
rect -212 -472 -206 -438
rect -252 -510 -206 -472
rect -252 -544 -246 -510
rect -212 -544 -206 -510
rect -252 -582 -206 -544
rect -252 -616 -246 -582
rect -212 -616 -206 -582
rect -252 -647 -206 -616
rect 206 -78 252 -47
rect 206 -112 212 -78
rect 246 -112 252 -78
rect 206 -150 252 -112
rect 206 -184 212 -150
rect 246 -184 252 -150
rect 206 -222 252 -184
rect 206 -256 212 -222
rect 246 -256 252 -222
rect 206 -294 252 -256
rect 206 -328 212 -294
rect 246 -328 252 -294
rect 206 -366 252 -328
rect 206 -400 212 -366
rect 246 -400 252 -366
rect 206 -438 252 -400
rect 206 -472 212 -438
rect 246 -472 252 -438
rect 206 -510 252 -472
rect 206 -544 212 -510
rect 246 -544 252 -510
rect 206 -582 252 -544
rect 206 -616 212 -582
rect 246 -616 252 -582
rect 206 -647 252 -616
rect 664 -78 710 -47
rect 664 -112 670 -78
rect 704 -112 710 -78
rect 664 -150 710 -112
rect 664 -184 670 -150
rect 704 -184 710 -150
rect 664 -222 710 -184
rect 664 -256 670 -222
rect 704 -256 710 -222
rect 664 -294 710 -256
rect 664 -328 670 -294
rect 704 -328 710 -294
rect 664 -366 710 -328
rect 664 -400 670 -366
rect 704 -400 710 -366
rect 664 -438 710 -400
rect 664 -472 670 -438
rect 704 -472 710 -438
rect 664 -510 710 -472
rect 664 -544 670 -510
rect 704 -544 710 -510
rect 664 -582 710 -544
rect 664 -616 670 -582
rect 704 -616 710 -582
rect 664 -647 710 -616
rect 1122 -78 1168 -47
rect 1122 -112 1128 -78
rect 1162 -112 1168 -78
rect 1122 -150 1168 -112
rect 1122 -184 1128 -150
rect 1162 -184 1168 -150
rect 1122 -222 1168 -184
rect 1122 -256 1128 -222
rect 1162 -256 1168 -222
rect 1122 -294 1168 -256
rect 1122 -328 1128 -294
rect 1162 -328 1168 -294
rect 1122 -366 1168 -328
rect 1122 -400 1128 -366
rect 1162 -400 1168 -366
rect 1122 -438 1168 -400
rect 1122 -472 1128 -438
rect 1162 -472 1168 -438
rect 1122 -510 1168 -472
rect 1122 -544 1128 -510
rect 1162 -544 1168 -510
rect 1122 -582 1168 -544
rect 1122 -616 1128 -582
rect 1162 -616 1168 -582
rect 1122 -647 1168 -616
rect -1112 -685 -720 -679
rect -1112 -719 -1077 -685
rect -1043 -719 -1005 -685
rect -971 -719 -933 -685
rect -899 -719 -861 -685
rect -827 -719 -789 -685
rect -755 -719 -720 -685
rect -1112 -725 -720 -719
rect -654 -685 -262 -679
rect -654 -719 -619 -685
rect -585 -719 -547 -685
rect -513 -719 -475 -685
rect -441 -719 -403 -685
rect -369 -719 -331 -685
rect -297 -719 -262 -685
rect -654 -725 -262 -719
rect -196 -685 196 -679
rect -196 -719 -161 -685
rect -127 -719 -89 -685
rect -55 -719 -17 -685
rect 17 -719 55 -685
rect 89 -719 127 -685
rect 161 -719 196 -685
rect -196 -725 196 -719
rect 262 -685 654 -679
rect 262 -719 297 -685
rect 331 -719 369 -685
rect 403 -719 441 -685
rect 475 -719 513 -685
rect 547 -719 585 -685
rect 619 -719 654 -685
rect 262 -725 654 -719
rect 720 -685 1112 -679
rect 720 -719 755 -685
rect 789 -719 827 -685
rect 861 -719 899 -685
rect 933 -719 971 -685
rect 1005 -719 1043 -685
rect 1077 -719 1112 -685
rect 720 -725 1112 -719
rect -1168 -834 -1122 -803
rect -1168 -868 -1162 -834
rect -1128 -868 -1122 -834
rect -1168 -906 -1122 -868
rect -1168 -940 -1162 -906
rect -1128 -940 -1122 -906
rect -1168 -978 -1122 -940
rect -1168 -1012 -1162 -978
rect -1128 -1012 -1122 -978
rect -1168 -1050 -1122 -1012
rect -1168 -1084 -1162 -1050
rect -1128 -1084 -1122 -1050
rect -1168 -1122 -1122 -1084
rect -1168 -1156 -1162 -1122
rect -1128 -1156 -1122 -1122
rect -1168 -1194 -1122 -1156
rect -1168 -1228 -1162 -1194
rect -1128 -1228 -1122 -1194
rect -1168 -1266 -1122 -1228
rect -1168 -1300 -1162 -1266
rect -1128 -1300 -1122 -1266
rect -1168 -1338 -1122 -1300
rect -1168 -1372 -1162 -1338
rect -1128 -1372 -1122 -1338
rect -1168 -1403 -1122 -1372
rect -710 -834 -664 -803
rect -710 -868 -704 -834
rect -670 -868 -664 -834
rect -710 -906 -664 -868
rect -710 -940 -704 -906
rect -670 -940 -664 -906
rect -710 -978 -664 -940
rect -710 -1012 -704 -978
rect -670 -1012 -664 -978
rect -710 -1050 -664 -1012
rect -710 -1084 -704 -1050
rect -670 -1084 -664 -1050
rect -710 -1122 -664 -1084
rect -710 -1156 -704 -1122
rect -670 -1156 -664 -1122
rect -710 -1194 -664 -1156
rect -710 -1228 -704 -1194
rect -670 -1228 -664 -1194
rect -710 -1266 -664 -1228
rect -710 -1300 -704 -1266
rect -670 -1300 -664 -1266
rect -710 -1338 -664 -1300
rect -710 -1372 -704 -1338
rect -670 -1372 -664 -1338
rect -710 -1403 -664 -1372
rect -252 -834 -206 -803
rect -252 -868 -246 -834
rect -212 -868 -206 -834
rect -252 -906 -206 -868
rect -252 -940 -246 -906
rect -212 -940 -206 -906
rect -252 -978 -206 -940
rect -252 -1012 -246 -978
rect -212 -1012 -206 -978
rect -252 -1050 -206 -1012
rect -252 -1084 -246 -1050
rect -212 -1084 -206 -1050
rect -252 -1122 -206 -1084
rect -252 -1156 -246 -1122
rect -212 -1156 -206 -1122
rect -252 -1194 -206 -1156
rect -252 -1228 -246 -1194
rect -212 -1228 -206 -1194
rect -252 -1266 -206 -1228
rect -252 -1300 -246 -1266
rect -212 -1300 -206 -1266
rect -252 -1338 -206 -1300
rect -252 -1372 -246 -1338
rect -212 -1372 -206 -1338
rect -252 -1403 -206 -1372
rect 206 -834 252 -803
rect 206 -868 212 -834
rect 246 -868 252 -834
rect 206 -906 252 -868
rect 206 -940 212 -906
rect 246 -940 252 -906
rect 206 -978 252 -940
rect 206 -1012 212 -978
rect 246 -1012 252 -978
rect 206 -1050 252 -1012
rect 206 -1084 212 -1050
rect 246 -1084 252 -1050
rect 206 -1122 252 -1084
rect 206 -1156 212 -1122
rect 246 -1156 252 -1122
rect 206 -1194 252 -1156
rect 206 -1228 212 -1194
rect 246 -1228 252 -1194
rect 206 -1266 252 -1228
rect 206 -1300 212 -1266
rect 246 -1300 252 -1266
rect 206 -1338 252 -1300
rect 206 -1372 212 -1338
rect 246 -1372 252 -1338
rect 206 -1403 252 -1372
rect 664 -834 710 -803
rect 664 -868 670 -834
rect 704 -868 710 -834
rect 664 -906 710 -868
rect 664 -940 670 -906
rect 704 -940 710 -906
rect 664 -978 710 -940
rect 664 -1012 670 -978
rect 704 -1012 710 -978
rect 664 -1050 710 -1012
rect 664 -1084 670 -1050
rect 704 -1084 710 -1050
rect 664 -1122 710 -1084
rect 664 -1156 670 -1122
rect 704 -1156 710 -1122
rect 664 -1194 710 -1156
rect 664 -1228 670 -1194
rect 704 -1228 710 -1194
rect 664 -1266 710 -1228
rect 664 -1300 670 -1266
rect 704 -1300 710 -1266
rect 664 -1338 710 -1300
rect 664 -1372 670 -1338
rect 704 -1372 710 -1338
rect 664 -1403 710 -1372
rect 1122 -834 1168 -803
rect 1122 -868 1128 -834
rect 1162 -868 1168 -834
rect 1122 -906 1168 -868
rect 1122 -940 1128 -906
rect 1162 -940 1168 -906
rect 1122 -978 1168 -940
rect 1122 -1012 1128 -978
rect 1162 -1012 1168 -978
rect 1122 -1050 1168 -1012
rect 1122 -1084 1128 -1050
rect 1162 -1084 1168 -1050
rect 1122 -1122 1168 -1084
rect 1122 -1156 1128 -1122
rect 1162 -1156 1168 -1122
rect 1122 -1194 1168 -1156
rect 1122 -1228 1128 -1194
rect 1162 -1228 1168 -1194
rect 1122 -1266 1168 -1228
rect 1122 -1300 1128 -1266
rect 1162 -1300 1168 -1266
rect 1122 -1338 1168 -1300
rect 1122 -1372 1128 -1338
rect 1162 -1372 1168 -1338
rect 1122 -1403 1168 -1372
rect -1112 -1441 -720 -1435
rect -1112 -1475 -1077 -1441
rect -1043 -1475 -1005 -1441
rect -971 -1475 -933 -1441
rect -899 -1475 -861 -1441
rect -827 -1475 -789 -1441
rect -755 -1475 -720 -1441
rect -1112 -1481 -720 -1475
rect -654 -1441 -262 -1435
rect -654 -1475 -619 -1441
rect -585 -1475 -547 -1441
rect -513 -1475 -475 -1441
rect -441 -1475 -403 -1441
rect -369 -1475 -331 -1441
rect -297 -1475 -262 -1441
rect -654 -1481 -262 -1475
rect -196 -1441 196 -1435
rect -196 -1475 -161 -1441
rect -127 -1475 -89 -1441
rect -55 -1475 -17 -1441
rect 17 -1475 55 -1441
rect 89 -1475 127 -1441
rect 161 -1475 196 -1441
rect -196 -1481 196 -1475
rect 262 -1441 654 -1435
rect 262 -1475 297 -1441
rect 331 -1475 369 -1441
rect 403 -1475 441 -1441
rect 475 -1475 513 -1441
rect 547 -1475 585 -1441
rect 619 -1475 654 -1441
rect 262 -1481 654 -1475
rect 720 -1441 1112 -1435
rect 720 -1475 755 -1441
rect 789 -1475 827 -1441
rect 861 -1475 899 -1441
rect 933 -1475 971 -1441
rect 1005 -1475 1043 -1441
rect 1077 -1475 1112 -1441
rect 720 -1481 1112 -1475
<< properties >>
string FIXED_BBOX -1259 -1560 1259 1560
<< end >>
