magic
tech sky130A
timestamp 1666387681
<< locali >>
rect 20 4410 3200 4440
rect 20 3960 3200 3990
rect 20 3770 3200 3800
rect 30 3310 3210 3340
rect 30 3120 3210 3150
rect 30 2670 3210 2700
rect 30 2480 3210 2510
rect 30 2030 3210 2060
rect 30 1830 3210 1860
rect 30 1380 3210 1410
rect 40 1190 3220 1220
rect 40 740 3220 770
rect 40 550 3220 580
rect 40 90 3220 120
<< metal1 >>
rect 300 4150 3000 4250
rect 600 3600 700 4150
rect 1250 3600 1350 4150
rect 1900 3600 2000 4150
rect 2550 3600 2650 4150
rect 300 3500 3000 3600
rect 600 2950 700 3500
rect 1250 2950 1350 3500
rect 1900 2950 2000 3500
rect 2550 2950 2650 3500
rect 300 2850 3000 2950
rect 600 2300 700 2850
rect 250 2200 1050 2300
rect 600 1650 700 2200
rect 1250 1650 1350 2850
rect 1545 2200 1550 2350
rect 1700 2200 1705 2350
rect 1900 1650 2000 2850
rect 2550 2300 2650 2850
rect 2200 2200 3000 2300
rect 2550 1650 2650 2200
rect 300 1550 3000 1650
rect 600 1000 700 1550
rect 1250 1000 1350 1550
rect 1900 1000 2000 1550
rect 2550 1000 2650 1550
rect 300 900 3000 1000
rect 600 400 700 900
rect 1250 400 1350 900
rect 1900 400 2000 900
rect 2550 400 2650 900
rect 250 300 2950 400
<< via1 >>
rect 1550 2200 1700 2350
<< metal2 >>
rect 1550 2350 1700 2355
rect 1550 2195 1700 2200
use sky130_fd_pr__rf_pnp_05v5_W3p40L3p40  sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0 $PDKPATH/libs.ref/sky130_fd_pr/mag
array 0 4 644 0 6 644
timestamp 1666199351
transform 1 0 0 0 1 0
box 0 0 670 670
<< end >>
