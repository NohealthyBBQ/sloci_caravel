magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< pwell >>
rect -571 -445 571 507
<< nmoslvt >>
rect -487 -419 -287 481
rect -229 -419 -29 481
rect 29 -419 229 481
rect 287 -419 487 481
<< ndiff >>
rect -545 456 -487 481
rect -545 422 -533 456
rect -499 422 -487 456
rect -545 388 -487 422
rect -545 354 -533 388
rect -499 354 -487 388
rect -545 320 -487 354
rect -545 286 -533 320
rect -499 286 -487 320
rect -545 252 -487 286
rect -545 218 -533 252
rect -499 218 -487 252
rect -545 184 -487 218
rect -545 150 -533 184
rect -499 150 -487 184
rect -545 116 -487 150
rect -545 82 -533 116
rect -499 82 -487 116
rect -545 48 -487 82
rect -545 14 -533 48
rect -499 14 -487 48
rect -545 -20 -487 14
rect -545 -54 -533 -20
rect -499 -54 -487 -20
rect -545 -88 -487 -54
rect -545 -122 -533 -88
rect -499 -122 -487 -88
rect -545 -156 -487 -122
rect -545 -190 -533 -156
rect -499 -190 -487 -156
rect -545 -224 -487 -190
rect -545 -258 -533 -224
rect -499 -258 -487 -224
rect -545 -292 -487 -258
rect -545 -326 -533 -292
rect -499 -326 -487 -292
rect -545 -360 -487 -326
rect -545 -394 -533 -360
rect -499 -394 -487 -360
rect -545 -419 -487 -394
rect -287 456 -229 481
rect -287 422 -275 456
rect -241 422 -229 456
rect -287 388 -229 422
rect -287 354 -275 388
rect -241 354 -229 388
rect -287 320 -229 354
rect -287 286 -275 320
rect -241 286 -229 320
rect -287 252 -229 286
rect -287 218 -275 252
rect -241 218 -229 252
rect -287 184 -229 218
rect -287 150 -275 184
rect -241 150 -229 184
rect -287 116 -229 150
rect -287 82 -275 116
rect -241 82 -229 116
rect -287 48 -229 82
rect -287 14 -275 48
rect -241 14 -229 48
rect -287 -20 -229 14
rect -287 -54 -275 -20
rect -241 -54 -229 -20
rect -287 -88 -229 -54
rect -287 -122 -275 -88
rect -241 -122 -229 -88
rect -287 -156 -229 -122
rect -287 -190 -275 -156
rect -241 -190 -229 -156
rect -287 -224 -229 -190
rect -287 -258 -275 -224
rect -241 -258 -229 -224
rect -287 -292 -229 -258
rect -287 -326 -275 -292
rect -241 -326 -229 -292
rect -287 -360 -229 -326
rect -287 -394 -275 -360
rect -241 -394 -229 -360
rect -287 -419 -229 -394
rect -29 456 29 481
rect -29 422 -17 456
rect 17 422 29 456
rect -29 388 29 422
rect -29 354 -17 388
rect 17 354 29 388
rect -29 320 29 354
rect -29 286 -17 320
rect 17 286 29 320
rect -29 252 29 286
rect -29 218 -17 252
rect 17 218 29 252
rect -29 184 29 218
rect -29 150 -17 184
rect 17 150 29 184
rect -29 116 29 150
rect -29 82 -17 116
rect 17 82 29 116
rect -29 48 29 82
rect -29 14 -17 48
rect 17 14 29 48
rect -29 -20 29 14
rect -29 -54 -17 -20
rect 17 -54 29 -20
rect -29 -88 29 -54
rect -29 -122 -17 -88
rect 17 -122 29 -88
rect -29 -156 29 -122
rect -29 -190 -17 -156
rect 17 -190 29 -156
rect -29 -224 29 -190
rect -29 -258 -17 -224
rect 17 -258 29 -224
rect -29 -292 29 -258
rect -29 -326 -17 -292
rect 17 -326 29 -292
rect -29 -360 29 -326
rect -29 -394 -17 -360
rect 17 -394 29 -360
rect -29 -419 29 -394
rect 229 456 287 481
rect 229 422 241 456
rect 275 422 287 456
rect 229 388 287 422
rect 229 354 241 388
rect 275 354 287 388
rect 229 320 287 354
rect 229 286 241 320
rect 275 286 287 320
rect 229 252 287 286
rect 229 218 241 252
rect 275 218 287 252
rect 229 184 287 218
rect 229 150 241 184
rect 275 150 287 184
rect 229 116 287 150
rect 229 82 241 116
rect 275 82 287 116
rect 229 48 287 82
rect 229 14 241 48
rect 275 14 287 48
rect 229 -20 287 14
rect 229 -54 241 -20
rect 275 -54 287 -20
rect 229 -88 287 -54
rect 229 -122 241 -88
rect 275 -122 287 -88
rect 229 -156 287 -122
rect 229 -190 241 -156
rect 275 -190 287 -156
rect 229 -224 287 -190
rect 229 -258 241 -224
rect 275 -258 287 -224
rect 229 -292 287 -258
rect 229 -326 241 -292
rect 275 -326 287 -292
rect 229 -360 287 -326
rect 229 -394 241 -360
rect 275 -394 287 -360
rect 229 -419 287 -394
rect 487 456 545 481
rect 487 422 499 456
rect 533 422 545 456
rect 487 388 545 422
rect 487 354 499 388
rect 533 354 545 388
rect 487 320 545 354
rect 487 286 499 320
rect 533 286 545 320
rect 487 252 545 286
rect 487 218 499 252
rect 533 218 545 252
rect 487 184 545 218
rect 487 150 499 184
rect 533 150 545 184
rect 487 116 545 150
rect 487 82 499 116
rect 533 82 545 116
rect 487 48 545 82
rect 487 14 499 48
rect 533 14 545 48
rect 487 -20 545 14
rect 487 -54 499 -20
rect 533 -54 545 -20
rect 487 -88 545 -54
rect 487 -122 499 -88
rect 533 -122 545 -88
rect 487 -156 545 -122
rect 487 -190 499 -156
rect 533 -190 545 -156
rect 487 -224 545 -190
rect 487 -258 499 -224
rect 533 -258 545 -224
rect 487 -292 545 -258
rect 487 -326 499 -292
rect 533 -326 545 -292
rect 487 -360 545 -326
rect 487 -394 499 -360
rect 533 -394 545 -360
rect 487 -419 545 -394
<< ndiffc >>
rect -533 422 -499 456
rect -533 354 -499 388
rect -533 286 -499 320
rect -533 218 -499 252
rect -533 150 -499 184
rect -533 82 -499 116
rect -533 14 -499 48
rect -533 -54 -499 -20
rect -533 -122 -499 -88
rect -533 -190 -499 -156
rect -533 -258 -499 -224
rect -533 -326 -499 -292
rect -533 -394 -499 -360
rect -275 422 -241 456
rect -275 354 -241 388
rect -275 286 -241 320
rect -275 218 -241 252
rect -275 150 -241 184
rect -275 82 -241 116
rect -275 14 -241 48
rect -275 -54 -241 -20
rect -275 -122 -241 -88
rect -275 -190 -241 -156
rect -275 -258 -241 -224
rect -275 -326 -241 -292
rect -275 -394 -241 -360
rect -17 422 17 456
rect -17 354 17 388
rect -17 286 17 320
rect -17 218 17 252
rect -17 150 17 184
rect -17 82 17 116
rect -17 14 17 48
rect -17 -54 17 -20
rect -17 -122 17 -88
rect -17 -190 17 -156
rect -17 -258 17 -224
rect -17 -326 17 -292
rect -17 -394 17 -360
rect 241 422 275 456
rect 241 354 275 388
rect 241 286 275 320
rect 241 218 275 252
rect 241 150 275 184
rect 241 82 275 116
rect 241 14 275 48
rect 241 -54 275 -20
rect 241 -122 275 -88
rect 241 -190 275 -156
rect 241 -258 275 -224
rect 241 -326 275 -292
rect 241 -394 275 -360
rect 499 422 533 456
rect 499 354 533 388
rect 499 286 533 320
rect 499 218 533 252
rect 499 150 533 184
rect 499 82 533 116
rect 499 14 533 48
rect 499 -54 533 -20
rect 499 -122 533 -88
rect 499 -190 533 -156
rect 499 -258 533 -224
rect 499 -326 533 -292
rect 499 -394 533 -360
<< poly >>
rect -487 481 -287 507
rect -229 481 -29 507
rect 29 481 229 507
rect 287 481 487 507
rect -487 -457 -287 -419
rect -487 -491 -438 -457
rect -404 -491 -370 -457
rect -336 -491 -287 -457
rect -487 -507 -287 -491
rect -229 -457 -29 -419
rect -229 -491 -180 -457
rect -146 -491 -112 -457
rect -78 -491 -29 -457
rect -229 -507 -29 -491
rect 29 -457 229 -419
rect 29 -491 78 -457
rect 112 -491 146 -457
rect 180 -491 229 -457
rect 29 -507 229 -491
rect 287 -457 487 -419
rect 287 -491 336 -457
rect 370 -491 404 -457
rect 438 -491 487 -457
rect 287 -507 487 -491
<< polycont >>
rect -438 -491 -404 -457
rect -370 -491 -336 -457
rect -180 -491 -146 -457
rect -112 -491 -78 -457
rect 78 -491 112 -457
rect 146 -491 180 -457
rect 336 -491 370 -457
rect 404 -491 438 -457
<< locali >>
rect -533 456 -499 485
rect -533 388 -499 410
rect -533 320 -499 338
rect -533 252 -499 266
rect -533 184 -499 194
rect -533 116 -499 122
rect -533 48 -499 50
rect -533 12 -499 14
rect -533 -60 -499 -54
rect -533 -132 -499 -122
rect -533 -204 -499 -190
rect -533 -276 -499 -258
rect -533 -348 -499 -326
rect -533 -423 -499 -394
rect -275 456 -241 485
rect -275 388 -241 410
rect -275 320 -241 338
rect -275 252 -241 266
rect -275 184 -241 194
rect -275 116 -241 122
rect -275 48 -241 50
rect -275 12 -241 14
rect -275 -60 -241 -54
rect -275 -132 -241 -122
rect -275 -204 -241 -190
rect -275 -276 -241 -258
rect -275 -348 -241 -326
rect -275 -423 -241 -394
rect -17 456 17 485
rect -17 388 17 410
rect -17 320 17 338
rect -17 252 17 266
rect -17 184 17 194
rect -17 116 17 122
rect -17 48 17 50
rect -17 12 17 14
rect -17 -60 17 -54
rect -17 -132 17 -122
rect -17 -204 17 -190
rect -17 -276 17 -258
rect -17 -348 17 -326
rect -17 -423 17 -394
rect 241 456 275 485
rect 241 388 275 410
rect 241 320 275 338
rect 241 252 275 266
rect 241 184 275 194
rect 241 116 275 122
rect 241 48 275 50
rect 241 12 275 14
rect 241 -60 275 -54
rect 241 -132 275 -122
rect 241 -204 275 -190
rect 241 -276 275 -258
rect 241 -348 275 -326
rect 241 -423 275 -394
rect 499 456 533 485
rect 499 388 533 410
rect 499 320 533 338
rect 499 252 533 266
rect 499 184 533 194
rect 499 116 533 122
rect 499 48 533 50
rect 499 12 533 14
rect 499 -60 533 -54
rect 499 -132 533 -122
rect 499 -204 533 -190
rect 499 -276 533 -258
rect 499 -348 533 -326
rect 499 -423 533 -394
rect -487 -491 -440 -457
rect -404 -491 -370 -457
rect -334 -491 -287 -457
rect -229 -491 -182 -457
rect -146 -491 -112 -457
rect -76 -491 -29 -457
rect 29 -491 76 -457
rect 112 -491 146 -457
rect 182 -491 229 -457
rect 287 -491 334 -457
rect 370 -491 404 -457
rect 440 -491 487 -457
<< viali >>
rect -533 422 -499 444
rect -533 410 -499 422
rect -533 354 -499 372
rect -533 338 -499 354
rect -533 286 -499 300
rect -533 266 -499 286
rect -533 218 -499 228
rect -533 194 -499 218
rect -533 150 -499 156
rect -533 122 -499 150
rect -533 82 -499 84
rect -533 50 -499 82
rect -533 -20 -499 12
rect -533 -22 -499 -20
rect -533 -88 -499 -60
rect -533 -94 -499 -88
rect -533 -156 -499 -132
rect -533 -166 -499 -156
rect -533 -224 -499 -204
rect -533 -238 -499 -224
rect -533 -292 -499 -276
rect -533 -310 -499 -292
rect -533 -360 -499 -348
rect -533 -382 -499 -360
rect -275 422 -241 444
rect -275 410 -241 422
rect -275 354 -241 372
rect -275 338 -241 354
rect -275 286 -241 300
rect -275 266 -241 286
rect -275 218 -241 228
rect -275 194 -241 218
rect -275 150 -241 156
rect -275 122 -241 150
rect -275 82 -241 84
rect -275 50 -241 82
rect -275 -20 -241 12
rect -275 -22 -241 -20
rect -275 -88 -241 -60
rect -275 -94 -241 -88
rect -275 -156 -241 -132
rect -275 -166 -241 -156
rect -275 -224 -241 -204
rect -275 -238 -241 -224
rect -275 -292 -241 -276
rect -275 -310 -241 -292
rect -275 -360 -241 -348
rect -275 -382 -241 -360
rect -17 422 17 444
rect -17 410 17 422
rect -17 354 17 372
rect -17 338 17 354
rect -17 286 17 300
rect -17 266 17 286
rect -17 218 17 228
rect -17 194 17 218
rect -17 150 17 156
rect -17 122 17 150
rect -17 82 17 84
rect -17 50 17 82
rect -17 -20 17 12
rect -17 -22 17 -20
rect -17 -88 17 -60
rect -17 -94 17 -88
rect -17 -156 17 -132
rect -17 -166 17 -156
rect -17 -224 17 -204
rect -17 -238 17 -224
rect -17 -292 17 -276
rect -17 -310 17 -292
rect -17 -360 17 -348
rect -17 -382 17 -360
rect 241 422 275 444
rect 241 410 275 422
rect 241 354 275 372
rect 241 338 275 354
rect 241 286 275 300
rect 241 266 275 286
rect 241 218 275 228
rect 241 194 275 218
rect 241 150 275 156
rect 241 122 275 150
rect 241 82 275 84
rect 241 50 275 82
rect 241 -20 275 12
rect 241 -22 275 -20
rect 241 -88 275 -60
rect 241 -94 275 -88
rect 241 -156 275 -132
rect 241 -166 275 -156
rect 241 -224 275 -204
rect 241 -238 275 -224
rect 241 -292 275 -276
rect 241 -310 275 -292
rect 241 -360 275 -348
rect 241 -382 275 -360
rect 499 422 533 444
rect 499 410 533 422
rect 499 354 533 372
rect 499 338 533 354
rect 499 286 533 300
rect 499 266 533 286
rect 499 218 533 228
rect 499 194 533 218
rect 499 150 533 156
rect 499 122 533 150
rect 499 82 533 84
rect 499 50 533 82
rect 499 -20 533 12
rect 499 -22 533 -20
rect 499 -88 533 -60
rect 499 -94 533 -88
rect 499 -156 533 -132
rect 499 -166 533 -156
rect 499 -224 533 -204
rect 499 -238 533 -224
rect 499 -292 533 -276
rect 499 -310 533 -292
rect 499 -360 533 -348
rect 499 -382 533 -360
rect -440 -491 -438 -457
rect -438 -491 -406 -457
rect -368 -491 -336 -457
rect -336 -491 -334 -457
rect -182 -491 -180 -457
rect -180 -491 -148 -457
rect -110 -491 -78 -457
rect -78 -491 -76 -457
rect 76 -491 78 -457
rect 78 -491 110 -457
rect 148 -491 180 -457
rect 180 -491 182 -457
rect 334 -491 336 -457
rect 336 -491 368 -457
rect 406 -491 438 -457
rect 438 -491 440 -457
<< metal1 >>
rect -539 444 -493 481
rect -539 410 -533 444
rect -499 410 -493 444
rect -539 372 -493 410
rect -539 338 -533 372
rect -499 338 -493 372
rect -539 300 -493 338
rect -539 266 -533 300
rect -499 266 -493 300
rect -539 228 -493 266
rect -539 194 -533 228
rect -499 194 -493 228
rect -539 156 -493 194
rect -539 122 -533 156
rect -499 122 -493 156
rect -539 84 -493 122
rect -539 50 -533 84
rect -499 50 -493 84
rect -539 12 -493 50
rect -539 -22 -533 12
rect -499 -22 -493 12
rect -539 -60 -493 -22
rect -539 -94 -533 -60
rect -499 -94 -493 -60
rect -539 -132 -493 -94
rect -539 -166 -533 -132
rect -499 -166 -493 -132
rect -539 -204 -493 -166
rect -539 -238 -533 -204
rect -499 -238 -493 -204
rect -539 -276 -493 -238
rect -539 -310 -533 -276
rect -499 -310 -493 -276
rect -539 -348 -493 -310
rect -539 -382 -533 -348
rect -499 -382 -493 -348
rect -539 -419 -493 -382
rect -281 444 -235 481
rect -281 410 -275 444
rect -241 410 -235 444
rect -281 372 -235 410
rect -281 338 -275 372
rect -241 338 -235 372
rect -281 300 -235 338
rect -281 266 -275 300
rect -241 266 -235 300
rect -281 228 -235 266
rect -281 194 -275 228
rect -241 194 -235 228
rect -281 156 -235 194
rect -281 122 -275 156
rect -241 122 -235 156
rect -281 84 -235 122
rect -281 50 -275 84
rect -241 50 -235 84
rect -281 12 -235 50
rect -281 -22 -275 12
rect -241 -22 -235 12
rect -281 -60 -235 -22
rect -281 -94 -275 -60
rect -241 -94 -235 -60
rect -281 -132 -235 -94
rect -281 -166 -275 -132
rect -241 -166 -235 -132
rect -281 -204 -235 -166
rect -281 -238 -275 -204
rect -241 -238 -235 -204
rect -281 -276 -235 -238
rect -281 -310 -275 -276
rect -241 -310 -235 -276
rect -281 -348 -235 -310
rect -281 -382 -275 -348
rect -241 -382 -235 -348
rect -281 -419 -235 -382
rect -23 444 23 481
rect -23 410 -17 444
rect 17 410 23 444
rect -23 372 23 410
rect -23 338 -17 372
rect 17 338 23 372
rect -23 300 23 338
rect -23 266 -17 300
rect 17 266 23 300
rect -23 228 23 266
rect -23 194 -17 228
rect 17 194 23 228
rect -23 156 23 194
rect -23 122 -17 156
rect 17 122 23 156
rect -23 84 23 122
rect -23 50 -17 84
rect 17 50 23 84
rect -23 12 23 50
rect -23 -22 -17 12
rect 17 -22 23 12
rect -23 -60 23 -22
rect -23 -94 -17 -60
rect 17 -94 23 -60
rect -23 -132 23 -94
rect -23 -166 -17 -132
rect 17 -166 23 -132
rect -23 -204 23 -166
rect -23 -238 -17 -204
rect 17 -238 23 -204
rect -23 -276 23 -238
rect -23 -310 -17 -276
rect 17 -310 23 -276
rect -23 -348 23 -310
rect -23 -382 -17 -348
rect 17 -382 23 -348
rect -23 -419 23 -382
rect 235 444 281 481
rect 235 410 241 444
rect 275 410 281 444
rect 235 372 281 410
rect 235 338 241 372
rect 275 338 281 372
rect 235 300 281 338
rect 235 266 241 300
rect 275 266 281 300
rect 235 228 281 266
rect 235 194 241 228
rect 275 194 281 228
rect 235 156 281 194
rect 235 122 241 156
rect 275 122 281 156
rect 235 84 281 122
rect 235 50 241 84
rect 275 50 281 84
rect 235 12 281 50
rect 235 -22 241 12
rect 275 -22 281 12
rect 235 -60 281 -22
rect 235 -94 241 -60
rect 275 -94 281 -60
rect 235 -132 281 -94
rect 235 -166 241 -132
rect 275 -166 281 -132
rect 235 -204 281 -166
rect 235 -238 241 -204
rect 275 -238 281 -204
rect 235 -276 281 -238
rect 235 -310 241 -276
rect 275 -310 281 -276
rect 235 -348 281 -310
rect 235 -382 241 -348
rect 275 -382 281 -348
rect 235 -419 281 -382
rect 493 444 539 481
rect 493 410 499 444
rect 533 410 539 444
rect 493 372 539 410
rect 493 338 499 372
rect 533 338 539 372
rect 493 300 539 338
rect 493 266 499 300
rect 533 266 539 300
rect 493 228 539 266
rect 493 194 499 228
rect 533 194 539 228
rect 493 156 539 194
rect 493 122 499 156
rect 533 122 539 156
rect 493 84 539 122
rect 493 50 499 84
rect 533 50 539 84
rect 493 12 539 50
rect 493 -22 499 12
rect 533 -22 539 12
rect 493 -60 539 -22
rect 493 -94 499 -60
rect 533 -94 539 -60
rect 493 -132 539 -94
rect 493 -166 499 -132
rect 533 -166 539 -132
rect 493 -204 539 -166
rect 493 -238 499 -204
rect 533 -238 539 -204
rect 493 -276 539 -238
rect 493 -310 499 -276
rect 533 -310 539 -276
rect 493 -348 539 -310
rect 493 -382 499 -348
rect 533 -382 539 -348
rect 493 -419 539 -382
rect -483 -457 -291 -451
rect -483 -491 -440 -457
rect -406 -491 -368 -457
rect -334 -491 -291 -457
rect -483 -497 -291 -491
rect -225 -457 -33 -451
rect -225 -491 -182 -457
rect -148 -491 -110 -457
rect -76 -491 -33 -457
rect -225 -497 -33 -491
rect 33 -457 225 -451
rect 33 -491 76 -457
rect 110 -491 148 -457
rect 182 -491 225 -457
rect 33 -497 225 -491
rect 291 -457 483 -451
rect 291 -491 334 -457
rect 368 -491 406 -457
rect 440 -491 483 -457
rect 291 -497 483 -491
<< end >>
