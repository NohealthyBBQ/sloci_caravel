magic
tech sky130A
magscale 1 2
timestamp 1663011646
<< error_p >>
rect -607 181 -545 187
rect -479 181 -417 187
rect -351 181 -289 187
rect -223 181 -161 187
rect -95 181 -33 187
rect 33 181 95 187
rect 161 181 223 187
rect 289 181 351 187
rect 417 181 479 187
rect 545 181 607 187
rect -607 147 -593 181
rect -479 147 -465 181
rect -351 147 -337 181
rect -223 147 -209 181
rect -95 147 -81 181
rect 33 147 47 181
rect 161 147 175 181
rect 289 147 303 181
rect 417 147 431 181
rect 545 147 559 181
rect -607 141 -545 147
rect -479 141 -417 147
rect -351 141 -289 147
rect -223 141 -161 147
rect -95 141 -33 147
rect 33 141 95 147
rect 161 141 223 147
rect 289 141 351 147
rect 417 141 479 147
rect 545 141 607 147
rect -607 -147 -545 -141
rect -479 -147 -417 -141
rect -351 -147 -289 -141
rect -223 -147 -161 -141
rect -95 -147 -33 -141
rect 33 -147 95 -141
rect 161 -147 223 -141
rect 289 -147 351 -141
rect 417 -147 479 -141
rect 545 -147 607 -141
rect -607 -181 -593 -147
rect -479 -181 -465 -147
rect -351 -181 -337 -147
rect -223 -181 -209 -147
rect -95 -181 -81 -147
rect 33 -181 47 -147
rect 161 -181 175 -147
rect 289 -181 303 -147
rect 417 -181 431 -147
rect 545 -181 559 -147
rect -607 -187 -545 -181
rect -479 -187 -417 -181
rect -351 -187 -289 -181
rect -223 -187 -161 -181
rect -95 -187 -33 -181
rect 33 -187 95 -181
rect 161 -187 223 -181
rect 289 -187 351 -181
rect 417 -187 479 -181
rect 545 -187 607 -181
<< nwell >>
rect -807 -319 807 319
<< pmoslvt >>
rect -611 -100 -541 100
rect -483 -100 -413 100
rect -355 -100 -285 100
rect -227 -100 -157 100
rect -99 -100 -29 100
rect 29 -100 99 100
rect 157 -100 227 100
rect 285 -100 355 100
rect 413 -100 483 100
rect 541 -100 611 100
<< pdiff >>
rect -669 85 -611 100
rect -669 51 -657 85
rect -623 51 -611 85
rect -669 17 -611 51
rect -669 -17 -657 17
rect -623 -17 -611 17
rect -669 -51 -611 -17
rect -669 -85 -657 -51
rect -623 -85 -611 -51
rect -669 -100 -611 -85
rect -541 85 -483 100
rect -541 51 -529 85
rect -495 51 -483 85
rect -541 17 -483 51
rect -541 -17 -529 17
rect -495 -17 -483 17
rect -541 -51 -483 -17
rect -541 -85 -529 -51
rect -495 -85 -483 -51
rect -541 -100 -483 -85
rect -413 85 -355 100
rect -413 51 -401 85
rect -367 51 -355 85
rect -413 17 -355 51
rect -413 -17 -401 17
rect -367 -17 -355 17
rect -413 -51 -355 -17
rect -413 -85 -401 -51
rect -367 -85 -355 -51
rect -413 -100 -355 -85
rect -285 85 -227 100
rect -285 51 -273 85
rect -239 51 -227 85
rect -285 17 -227 51
rect -285 -17 -273 17
rect -239 -17 -227 17
rect -285 -51 -227 -17
rect -285 -85 -273 -51
rect -239 -85 -227 -51
rect -285 -100 -227 -85
rect -157 85 -99 100
rect -157 51 -145 85
rect -111 51 -99 85
rect -157 17 -99 51
rect -157 -17 -145 17
rect -111 -17 -99 17
rect -157 -51 -99 -17
rect -157 -85 -145 -51
rect -111 -85 -99 -51
rect -157 -100 -99 -85
rect -29 85 29 100
rect -29 51 -17 85
rect 17 51 29 85
rect -29 17 29 51
rect -29 -17 -17 17
rect 17 -17 29 17
rect -29 -51 29 -17
rect -29 -85 -17 -51
rect 17 -85 29 -51
rect -29 -100 29 -85
rect 99 85 157 100
rect 99 51 111 85
rect 145 51 157 85
rect 99 17 157 51
rect 99 -17 111 17
rect 145 -17 157 17
rect 99 -51 157 -17
rect 99 -85 111 -51
rect 145 -85 157 -51
rect 99 -100 157 -85
rect 227 85 285 100
rect 227 51 239 85
rect 273 51 285 85
rect 227 17 285 51
rect 227 -17 239 17
rect 273 -17 285 17
rect 227 -51 285 -17
rect 227 -85 239 -51
rect 273 -85 285 -51
rect 227 -100 285 -85
rect 355 85 413 100
rect 355 51 367 85
rect 401 51 413 85
rect 355 17 413 51
rect 355 -17 367 17
rect 401 -17 413 17
rect 355 -51 413 -17
rect 355 -85 367 -51
rect 401 -85 413 -51
rect 355 -100 413 -85
rect 483 85 541 100
rect 483 51 495 85
rect 529 51 541 85
rect 483 17 541 51
rect 483 -17 495 17
rect 529 -17 541 17
rect 483 -51 541 -17
rect 483 -85 495 -51
rect 529 -85 541 -51
rect 483 -100 541 -85
rect 611 85 669 100
rect 611 51 623 85
rect 657 51 669 85
rect 611 17 669 51
rect 611 -17 623 17
rect 657 -17 669 17
rect 611 -51 669 -17
rect 611 -85 623 -51
rect 657 -85 669 -51
rect 611 -100 669 -85
<< pdiffc >>
rect -657 51 -623 85
rect -657 -17 -623 17
rect -657 -85 -623 -51
rect -529 51 -495 85
rect -529 -17 -495 17
rect -529 -85 -495 -51
rect -401 51 -367 85
rect -401 -17 -367 17
rect -401 -85 -367 -51
rect -273 51 -239 85
rect -273 -17 -239 17
rect -273 -85 -239 -51
rect -145 51 -111 85
rect -145 -17 -111 17
rect -145 -85 -111 -51
rect -17 51 17 85
rect -17 -17 17 17
rect -17 -85 17 -51
rect 111 51 145 85
rect 111 -17 145 17
rect 111 -85 145 -51
rect 239 51 273 85
rect 239 -17 273 17
rect 239 -85 273 -51
rect 367 51 401 85
rect 367 -17 401 17
rect 367 -85 401 -51
rect 495 51 529 85
rect 495 -17 529 17
rect 495 -85 529 -51
rect 623 51 657 85
rect 623 -17 657 17
rect 623 -85 657 -51
<< nsubdiff >>
rect -771 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 771 283
rect -771 187 -737 249
rect -771 119 -737 153
rect 737 187 771 249
rect 737 119 771 153
rect -771 51 -737 85
rect -771 -17 -737 17
rect -771 -85 -737 -51
rect 737 51 771 85
rect 737 -17 771 17
rect 737 -85 771 -51
rect -771 -153 -737 -119
rect -771 -249 -737 -187
rect 737 -153 771 -119
rect 737 -249 771 -187
rect -771 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 771 -249
<< nsubdiffcont >>
rect -663 249 -629 283
rect -595 249 -561 283
rect -527 249 -493 283
rect -459 249 -425 283
rect -391 249 -357 283
rect -323 249 -289 283
rect -255 249 -221 283
rect -187 249 -153 283
rect -119 249 -85 283
rect -51 249 -17 283
rect 17 249 51 283
rect 85 249 119 283
rect 153 249 187 283
rect 221 249 255 283
rect 289 249 323 283
rect 357 249 391 283
rect 425 249 459 283
rect 493 249 527 283
rect 561 249 595 283
rect 629 249 663 283
rect -771 153 -737 187
rect -771 85 -737 119
rect 737 153 771 187
rect -771 17 -737 51
rect -771 -51 -737 -17
rect -771 -119 -737 -85
rect 737 85 771 119
rect 737 17 771 51
rect 737 -51 771 -17
rect -771 -187 -737 -153
rect 737 -119 771 -85
rect 737 -187 771 -153
rect -663 -283 -629 -249
rect -595 -283 -561 -249
rect -527 -283 -493 -249
rect -459 -283 -425 -249
rect -391 -283 -357 -249
rect -323 -283 -289 -249
rect -255 -283 -221 -249
rect -187 -283 -153 -249
rect -119 -283 -85 -249
rect -51 -283 -17 -249
rect 17 -283 51 -249
rect 85 -283 119 -249
rect 153 -283 187 -249
rect 221 -283 255 -249
rect 289 -283 323 -249
rect 357 -283 391 -249
rect 425 -283 459 -249
rect 493 -283 527 -249
rect 561 -283 595 -249
rect 629 -283 663 -249
<< poly >>
rect -611 181 -541 197
rect -611 147 -593 181
rect -559 147 -541 181
rect -611 100 -541 147
rect -483 181 -413 197
rect -483 147 -465 181
rect -431 147 -413 181
rect -483 100 -413 147
rect -355 181 -285 197
rect -355 147 -337 181
rect -303 147 -285 181
rect -355 100 -285 147
rect -227 181 -157 197
rect -227 147 -209 181
rect -175 147 -157 181
rect -227 100 -157 147
rect -99 181 -29 197
rect -99 147 -81 181
rect -47 147 -29 181
rect -99 100 -29 147
rect 29 181 99 197
rect 29 147 47 181
rect 81 147 99 181
rect 29 100 99 147
rect 157 181 227 197
rect 157 147 175 181
rect 209 147 227 181
rect 157 100 227 147
rect 285 181 355 197
rect 285 147 303 181
rect 337 147 355 181
rect 285 100 355 147
rect 413 181 483 197
rect 413 147 431 181
rect 465 147 483 181
rect 413 100 483 147
rect 541 181 611 197
rect 541 147 559 181
rect 593 147 611 181
rect 541 100 611 147
rect -611 -147 -541 -100
rect -611 -181 -593 -147
rect -559 -181 -541 -147
rect -611 -197 -541 -181
rect -483 -147 -413 -100
rect -483 -181 -465 -147
rect -431 -181 -413 -147
rect -483 -197 -413 -181
rect -355 -147 -285 -100
rect -355 -181 -337 -147
rect -303 -181 -285 -147
rect -355 -197 -285 -181
rect -227 -147 -157 -100
rect -227 -181 -209 -147
rect -175 -181 -157 -147
rect -227 -197 -157 -181
rect -99 -147 -29 -100
rect -99 -181 -81 -147
rect -47 -181 -29 -147
rect -99 -197 -29 -181
rect 29 -147 99 -100
rect 29 -181 47 -147
rect 81 -181 99 -147
rect 29 -197 99 -181
rect 157 -147 227 -100
rect 157 -181 175 -147
rect 209 -181 227 -147
rect 157 -197 227 -181
rect 285 -147 355 -100
rect 285 -181 303 -147
rect 337 -181 355 -147
rect 285 -197 355 -181
rect 413 -147 483 -100
rect 413 -181 431 -147
rect 465 -181 483 -147
rect 413 -197 483 -181
rect 541 -147 611 -100
rect 541 -181 559 -147
rect 593 -181 611 -147
rect 541 -197 611 -181
<< polycont >>
rect -593 147 -559 181
rect -465 147 -431 181
rect -337 147 -303 181
rect -209 147 -175 181
rect -81 147 -47 181
rect 47 147 81 181
rect 175 147 209 181
rect 303 147 337 181
rect 431 147 465 181
rect 559 147 593 181
rect -593 -181 -559 -147
rect -465 -181 -431 -147
rect -337 -181 -303 -147
rect -209 -181 -175 -147
rect -81 -181 -47 -147
rect 47 -181 81 -147
rect 175 -181 209 -147
rect 303 -181 337 -147
rect 431 -181 465 -147
rect 559 -181 593 -147
<< locali >>
rect -771 249 -663 283
rect -629 249 -595 283
rect -561 249 -527 283
rect -493 249 -459 283
rect -425 249 -391 283
rect -357 249 -323 283
rect -289 249 -255 283
rect -221 249 -187 283
rect -153 249 -119 283
rect -85 249 -51 283
rect -17 249 17 283
rect 51 249 85 283
rect 119 249 153 283
rect 187 249 221 283
rect 255 249 289 283
rect 323 249 357 283
rect 391 249 425 283
rect 459 249 493 283
rect 527 249 561 283
rect 595 249 629 283
rect 663 249 771 283
rect -771 187 -737 249
rect 737 187 771 249
rect -771 119 -737 153
rect -611 147 -593 181
rect -559 147 -541 181
rect -483 147 -465 181
rect -431 147 -413 181
rect -355 147 -337 181
rect -303 147 -285 181
rect -227 147 -209 181
rect -175 147 -157 181
rect -99 147 -81 181
rect -47 147 -29 181
rect 29 147 47 181
rect 81 147 99 181
rect 157 147 175 181
rect 209 147 227 181
rect 285 147 303 181
rect 337 147 355 181
rect 413 147 431 181
rect 465 147 483 181
rect 541 147 559 181
rect 593 147 611 181
rect 737 119 771 153
rect -771 51 -737 85
rect -771 -17 -737 17
rect -771 -85 -737 -51
rect -657 85 -623 104
rect -657 17 -623 19
rect -657 -19 -623 -17
rect -657 -104 -623 -85
rect -529 85 -495 104
rect -529 17 -495 19
rect -529 -19 -495 -17
rect -529 -104 -495 -85
rect -401 85 -367 104
rect -401 17 -367 19
rect -401 -19 -367 -17
rect -401 -104 -367 -85
rect -273 85 -239 104
rect -273 17 -239 19
rect -273 -19 -239 -17
rect -273 -104 -239 -85
rect -145 85 -111 104
rect -145 17 -111 19
rect -145 -19 -111 -17
rect -145 -104 -111 -85
rect -17 85 17 104
rect -17 17 17 19
rect -17 -19 17 -17
rect -17 -104 17 -85
rect 111 85 145 104
rect 111 17 145 19
rect 111 -19 145 -17
rect 111 -104 145 -85
rect 239 85 273 104
rect 239 17 273 19
rect 239 -19 273 -17
rect 239 -104 273 -85
rect 367 85 401 104
rect 367 17 401 19
rect 367 -19 401 -17
rect 367 -104 401 -85
rect 495 85 529 104
rect 495 17 529 19
rect 495 -19 529 -17
rect 495 -104 529 -85
rect 623 85 657 104
rect 623 17 657 19
rect 623 -19 657 -17
rect 623 -104 657 -85
rect 737 51 771 85
rect 737 -17 771 17
rect 737 -85 771 -51
rect -771 -153 -737 -119
rect -611 -181 -593 -147
rect -559 -181 -541 -147
rect -483 -181 -465 -147
rect -431 -181 -413 -147
rect -355 -181 -337 -147
rect -303 -181 -285 -147
rect -227 -181 -209 -147
rect -175 -181 -157 -147
rect -99 -181 -81 -147
rect -47 -181 -29 -147
rect 29 -181 47 -147
rect 81 -181 99 -147
rect 157 -181 175 -147
rect 209 -181 227 -147
rect 285 -181 303 -147
rect 337 -181 355 -147
rect 413 -181 431 -147
rect 465 -181 483 -147
rect 541 -181 559 -147
rect 593 -181 611 -147
rect 737 -153 771 -119
rect -771 -249 -737 -187
rect 737 -249 771 -187
rect -771 -283 -663 -249
rect -629 -283 -595 -249
rect -561 -283 -527 -249
rect -493 -283 -459 -249
rect -425 -283 -391 -249
rect -357 -283 -323 -249
rect -289 -283 -255 -249
rect -221 -283 -187 -249
rect -153 -283 -119 -249
rect -85 -283 -51 -249
rect -17 -283 17 -249
rect 51 -283 85 -249
rect 119 -283 153 -249
rect 187 -283 221 -249
rect 255 -283 289 -249
rect 323 -283 357 -249
rect 391 -283 425 -249
rect 459 -283 493 -249
rect 527 -283 561 -249
rect 595 -283 629 -249
rect 663 -283 771 -249
<< viali >>
rect -593 147 -559 181
rect -465 147 -431 181
rect -337 147 -303 181
rect -209 147 -175 181
rect -81 147 -47 181
rect 47 147 81 181
rect 175 147 209 181
rect 303 147 337 181
rect 431 147 465 181
rect 559 147 593 181
rect -657 51 -623 53
rect -657 19 -623 51
rect -657 -51 -623 -19
rect -657 -53 -623 -51
rect -529 51 -495 53
rect -529 19 -495 51
rect -529 -51 -495 -19
rect -529 -53 -495 -51
rect -401 51 -367 53
rect -401 19 -367 51
rect -401 -51 -367 -19
rect -401 -53 -367 -51
rect -273 51 -239 53
rect -273 19 -239 51
rect -273 -51 -239 -19
rect -273 -53 -239 -51
rect -145 51 -111 53
rect -145 19 -111 51
rect -145 -51 -111 -19
rect -145 -53 -111 -51
rect -17 51 17 53
rect -17 19 17 51
rect -17 -51 17 -19
rect -17 -53 17 -51
rect 111 51 145 53
rect 111 19 145 51
rect 111 -51 145 -19
rect 111 -53 145 -51
rect 239 51 273 53
rect 239 19 273 51
rect 239 -51 273 -19
rect 239 -53 273 -51
rect 367 51 401 53
rect 367 19 401 51
rect 367 -51 401 -19
rect 367 -53 401 -51
rect 495 51 529 53
rect 495 19 529 51
rect 495 -51 529 -19
rect 495 -53 529 -51
rect 623 51 657 53
rect 623 19 657 51
rect 623 -51 657 -19
rect 623 -53 657 -51
rect -593 -181 -559 -147
rect -465 -181 -431 -147
rect -337 -181 -303 -147
rect -209 -181 -175 -147
rect -81 -181 -47 -147
rect 47 -181 81 -147
rect 175 -181 209 -147
rect 303 -181 337 -147
rect 431 -181 465 -147
rect 559 -181 593 -147
<< metal1 >>
rect -607 181 -545 187
rect -607 147 -593 181
rect -559 147 -545 181
rect -607 141 -545 147
rect -479 181 -417 187
rect -479 147 -465 181
rect -431 147 -417 181
rect -479 141 -417 147
rect -351 181 -289 187
rect -351 147 -337 181
rect -303 147 -289 181
rect -351 141 -289 147
rect -223 181 -161 187
rect -223 147 -209 181
rect -175 147 -161 181
rect -223 141 -161 147
rect -95 181 -33 187
rect -95 147 -81 181
rect -47 147 -33 181
rect -95 141 -33 147
rect 33 181 95 187
rect 33 147 47 181
rect 81 147 95 181
rect 33 141 95 147
rect 161 181 223 187
rect 161 147 175 181
rect 209 147 223 181
rect 161 141 223 147
rect 289 181 351 187
rect 289 147 303 181
rect 337 147 351 181
rect 289 141 351 147
rect 417 181 479 187
rect 417 147 431 181
rect 465 147 479 181
rect 417 141 479 147
rect 545 181 607 187
rect 545 147 559 181
rect 593 147 607 181
rect 545 141 607 147
rect -663 53 -617 100
rect -663 19 -657 53
rect -623 19 -617 53
rect -663 -19 -617 19
rect -663 -53 -657 -19
rect -623 -53 -617 -19
rect -663 -100 -617 -53
rect -535 53 -489 100
rect -535 19 -529 53
rect -495 19 -489 53
rect -535 -19 -489 19
rect -535 -53 -529 -19
rect -495 -53 -489 -19
rect -535 -100 -489 -53
rect -407 53 -361 100
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -100 -361 -53
rect -279 53 -233 100
rect -279 19 -273 53
rect -239 19 -233 53
rect -279 -19 -233 19
rect -279 -53 -273 -19
rect -239 -53 -233 -19
rect -279 -100 -233 -53
rect -151 53 -105 100
rect -151 19 -145 53
rect -111 19 -105 53
rect -151 -19 -105 19
rect -151 -53 -145 -19
rect -111 -53 -105 -19
rect -151 -100 -105 -53
rect -23 53 23 100
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -100 23 -53
rect 105 53 151 100
rect 105 19 111 53
rect 145 19 151 53
rect 105 -19 151 19
rect 105 -53 111 -19
rect 145 -53 151 -19
rect 105 -100 151 -53
rect 233 53 279 100
rect 233 19 239 53
rect 273 19 279 53
rect 233 -19 279 19
rect 233 -53 239 -19
rect 273 -53 279 -19
rect 233 -100 279 -53
rect 361 53 407 100
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -100 407 -53
rect 489 53 535 100
rect 489 19 495 53
rect 529 19 535 53
rect 489 -19 535 19
rect 489 -53 495 -19
rect 529 -53 535 -19
rect 489 -100 535 -53
rect 617 53 663 100
rect 617 19 623 53
rect 657 19 663 53
rect 617 -19 663 19
rect 617 -53 623 -19
rect 657 -53 663 -19
rect 617 -100 663 -53
rect -607 -147 -545 -141
rect -607 -181 -593 -147
rect -559 -181 -545 -147
rect -607 -187 -545 -181
rect -479 -147 -417 -141
rect -479 -181 -465 -147
rect -431 -181 -417 -147
rect -479 -187 -417 -181
rect -351 -147 -289 -141
rect -351 -181 -337 -147
rect -303 -181 -289 -147
rect -351 -187 -289 -181
rect -223 -147 -161 -141
rect -223 -181 -209 -147
rect -175 -181 -161 -147
rect -223 -187 -161 -181
rect -95 -147 -33 -141
rect -95 -181 -81 -147
rect -47 -181 -33 -147
rect -95 -187 -33 -181
rect 33 -147 95 -141
rect 33 -181 47 -147
rect 81 -181 95 -147
rect 33 -187 95 -181
rect 161 -147 223 -141
rect 161 -181 175 -147
rect 209 -181 223 -147
rect 161 -187 223 -181
rect 289 -147 351 -141
rect 289 -181 303 -147
rect 337 -181 351 -147
rect 289 -187 351 -181
rect 417 -147 479 -141
rect 417 -181 431 -147
rect 465 -181 479 -147
rect 417 -187 479 -181
rect 545 -147 607 -141
rect 545 -181 559 -147
rect 593 -181 607 -147
rect 545 -187 607 -181
<< properties >>
string FIXED_BBOX -754 -266 754 266
<< end >>
